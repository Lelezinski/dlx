package alu_type is
  type alu_op_t is (ALU_ADD, ALU_SUB, ALU_AND, ALU_OR, ALU_XOR, ALU_SLL,
  ALU_SRL, ALU_SGE, ALU_SLE, ALU_SNE, ALU_MUL);
end alu_type;

-------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.constants.ALL;

-------------------------------------------------------------------------------

ENTITY ACC IS
	GENERIC (
		NBIT : INTEGER := numBit);
	PORT (
		A : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
		CLK : IN STD_LOGIC;
		RST_n : IN STD_LOGIC;
		ACCUMULATE : IN STD_LOGIC;
		ACC_EN_n : IN STD_LOGIC;
		Y : OUT STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0));
END ACC;

-------------------------------------------------------------------------------
-- Behavioral Architecture

ARCHITECTURE BEHAVIORAL OF ACC IS

	SIGNAL REG : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SIGNAL OUT_MUX : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SIGNAL OUT_ADD : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);

BEGIN
	MUX_PROCESS : PROCESS (B, REG, ACCUMULATE)
	BEGIN
		IF (ACCUMULATE = '1') THEN
			OUT_MUX <= REG;
		ELSE
			OUT_MUX <= B;
		END IF;
	END PROCESS;

	ADD_PROCESS : PROCESS (A, OUT_MUX)
	BEGIN
		OUT_ADD <= STD_LOGIC_VECTOR(unsigned(A) + unsigned(OUT_MUX));
	END PROCESS;

	REG_PROCESS : PROCESS (CLK, RST_n)
	BEGIN
		IF (RST_n = '0') THEN
			-- Async reset
			REG <= (OTHERS => '0');
		ELSIF (rising_edge(CLK)) THEN
			IF (ACC_EN_n = '0') THEN
				REG <= OUT_ADD;
			ELSE
				REG <= REG;
			END IF;
		END IF;
	END PROCESS;

	-- Output
	Y <= REG;

END BEHAVIORAL;

-------------------------------------------------------------------------------
-- Structural Architecture

ARCHITECTURE STRUCTURAL OF ACC IS

	SIGNAL FEED_BACK : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SIGNAL OUT_MUX : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SIGNAL OUT_ADD : STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SIGNAL RST : STD_LOGIC;

	-- Second Input MUX
	COMPONENT MUX21_GENERIC
		GENERIC (
			NBIT : INTEGER := numBit;
			DELAY_MUX : TIME := tp_mux);
		PORT (
			A : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			SEL : IN STD_LOGIC;
			Y : OUT STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0));
	END COMPONENT;

	-- Ripple Carry Adder
	COMPONENT RCA
		GENERIC (
			NBIT : INTEGER := numBit;
			DRCAS : TIME := 0 ns;
			DRCAC : TIME := 0 ns);
		PORT (
			A : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			Ci : IN STD_LOGIC;
			S : OUT STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			Co : OUT STD_LOGIC);
	END COMPONENT;

	-- Register Flip-Flop
	COMPONENT FD
		GENERIC (
			NBIT : INTEGER := numBit);
		PORT (
			D : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
			CK : IN STD_LOGIC;
			RESET : IN STD_LOGIC;
			Q : OUT STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0));
	END COMPONENT;

	-- Inverter (needed to match the active low reset)
	COMPONENT IV
		PORT (
			A : IN STD_LOGIC;
			Y : OUT STD_LOGIC);
	END COMPONENT;

BEGIN

	UMUX : MUX21_GENERIC
	PORT MAP(B, FEED_BACK, ACCUMULATE, OUT_MUX);

	URCA : RCA
	PORT MAP(A, OUT_MUX, '0', OUT_ADD, OPEN);

	UFD : FD
	PORT MAP(OUT_ADD, CLK, RST, FEED_BACK);

	UIV : IV
	PORT MAP(RST_n, RST);

	-- Output
	Y <= FEED_BACK;

END STRUCTURAL;

-------------------------------------------------------------------------------
-- Configs

CONFIGURATION CFG_ACC_BEHAVIORAL OF ACC IS
	FOR BEHAVIORAL
	END FOR;
END CFG_ACC_BEHAVIORAL;

CONFIGURATION CFG_ACC_STRUCTURAL OF ACC IS
	FOR STRUCTURAL
		FOR ALL : MUX21_GENERIC
		USE CONFIGURATION WORK.CFG_MUX21_GEN_STRUCTURAL;
	END FOR;
	FOR ALL : RCA
		USE CONFIGURATION WORK.CFG_RCA_STRUCTURAL;
	END FOR;
	FOR ALL : FD
		USE CONFIGURATION WORK.CFG_FD_PLUTO;
	END FOR;
	FOR ALL : IV
		USE CONFIGURATION WORK.CFG_IV_BEHAVIORAL;
	END FOR;
END FOR;
END CFG_ACC_STRUCTURAL;
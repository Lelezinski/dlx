
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_WINDOWED_REGISTER_FILE is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_WINDOWED_REGISTER_FILE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WINDOWED_REGISTER_FILE.all;

entity WINDOWED_REGISTER_FILE_DW01_addsub_0_DW01_addsub_2 is

   port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (4 downto 0);  CO : out std_logic);

end WINDOWED_REGISTER_FILE_DW01_addsub_0_DW01_addsub_2;

architecture SYN_rpl of WINDOWED_REGISTER_FILE_DW01_addsub_0_DW01_addsub_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_3_port, 
      B_AS_2_port, B_AS_1_port, B_AS_0_port, n_1003 : std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => ADD_SUB, CI => carry_4_port, CO => 
                           n_1003, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U2 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U3 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U4 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WINDOWED_REGISTER_FILE.all;

entity WINDOWED_REGISTER_FILE is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (3 downto 0);  DATAIN : in 
         std_logic_vector (7 downto 0);  OUT1, OUT2 : out std_logic_vector (7 
         downto 0);  CALL, RET : in std_logic;  FILL, SPILL : out std_logic;  
         FROM_MEM : in std_logic_vector (7 downto 0);  TO_MEM : out 
         std_logic_vector (7 downto 0));

end WINDOWED_REGISTER_FILE;

architecture SYN_BEHAVIORAL of WINDOWED_REGISTER_FILE is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component WINDOWED_REGISTER_FILE_DW01_addsub_0_DW01_addsub_2
      port( A, B : in std_logic_vector (4 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (4 downto 0);  CO : out 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal CWP_4_port, CWP_3_port, CWP_2_port, CWP_1_port, CWP_0_port, N201, 
      N202, N1662, N1663, N1664, N1665, N1666, n10, U3_U22_Z_0, U3_U22_Z_1, 
      U3_U22_Z_2, U3_U22_Z_3, U3_U23_Z_0, n1247, n1248, n1249, n1250, n1251, 
      n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, 
      n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, 
      n1272, n1273, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, 
      n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, 
      n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662_port, 
      n1663_port, n1664_port, n1665_port, n1666_port, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
      n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
      n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
      n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
      n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
      n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
      n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
      n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
      n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
      n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
      n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
      n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, 
      n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
      n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, 
      n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
      n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
      n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
      n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
      n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
      n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
      n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, 
      n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
      n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
      n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
      n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
      n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, 
      n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
      n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
      n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
      n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
      n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, 
      n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
      n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, 
      n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, 
      n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
      n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
      n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
      n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
      n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
      n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
      n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
      n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
      n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
      n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
      n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
      n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
      n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
      n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
      n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
      n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
      n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
      n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
      n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
      n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
      n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
      n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
      n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
      n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
      n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, SPILL_port, FILL_port, 
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094 : std_logic;

begin
   FILL <= FILL_port;
   SPILL <= SPILL_port;
   
   n10 <= '0';
   CANSAVE_reg_0_inst : DFF_X1 port map( D => n1797, CK => n2047, Q => n3285, 
                           QN => n_1004);
   STATE_reg_0_inst : DFF_X1 port map( D => N201, CK => n2050, Q => n3283, QN 
                           => n_1005);
   SWP_reg_0_inst : DFF_X1 port map( D => n1793, CK => n2047, Q => n1798, QN =>
                           n1495);
   STATE_reg_1_inst : DFF_X1 port map( D => N202, CK => n2047, Q => n3286, QN 
                           => n1944);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n1752, CK => n2047, Q => 
                           n_1006, QN => n1933);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n1753, CK => n2047, Q => 
                           n_1007, QN => n1924);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n1754, CK => n2047, Q => 
                           n_1008, QN => n1923);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n1755, CK => n2047, Q => 
                           n_1009, QN => n1922);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n1756, CK => n2048, Q => 
                           n_1010, QN => n1921);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n1757, CK => n2048, Q => 
                           n_1011, QN => n1920);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n1758, CK => n2048, Q => 
                           n_1012, QN => n1919);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n1759, CK => n2048, Q => 
                           n_1013, QN => n1918);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n1760, CK => n2048, Q => 
                           n3101, QN => n2035);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n1761, CK => n2048, Q => 
                           n3102, QN => n2042);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n1762, CK => n2048, Q => 
                           n3103, QN => n2041);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n1763, CK => n2048, Q => 
                           n3104, QN => n2040);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n1764, CK => n2048, Q => 
                           n3105, QN => n2039);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n1765, CK => n2048, Q => 
                           n3106, QN => n2038);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n1766, CK => n2048, Q => 
                           n3107, QN => n2037);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n1767, CK => n2049, Q => 
                           n3108, QN => n2036);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n1768, CK => n2049, Q => 
                           n_1014, QN => n3044);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n1769, CK => n2049, Q => 
                           n_1015, QN => n3043);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n1770, CK => n2049, Q => 
                           n_1016, QN => n3042);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n1771, CK => n2049, Q => 
                           n_1017, QN => n3041);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n1772, CK => n2049, Q => 
                           n_1018, QN => n3040);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n1773, CK => n2049, Q => 
                           n_1019, QN => n3039);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n1774, CK => n2049, Q => 
                           n_1020, QN => n3038);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n1775, CK => n2049, Q => 
                           n_1021, QN => n3037);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n1776, CK => n2049, Q => 
                           n1936, QN => n3219);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n1777, CK => n2049, Q => 
                           n1945, QN => n3225);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n1778, CK => n2050, Q => 
                           n1946, QN => n3233);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n1779, CK => n2050, Q => 
                           n1950, QN => n3241);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n1780, CK => n2050, Q => 
                           n1949, QN => n3249);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n1781, CK => n2050, Q => 
                           n1948, QN => n3257);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n1782, CK => n2050, Q => 
                           n1947, QN => n3265);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n1783, CK => n2050, Q => 
                           n1951, QN => n3273);
   CANRESTORE_reg_0_inst : DFF_X1 port map( D => n1795, CK => n2047, Q => n3281
                           , QN => n_1022);
   CANRESTORE_reg_1_inst : DFF_X1 port map( D => n1794, CK => n2047, Q => n3282
                           , QN => n_1023);
   SWP_reg_1_inst : DFF_X1 port map( D => n1792, CK => n2047, Q => n1830, QN =>
                           n1494);
   SWP_reg_4_inst : DFF_X1 port map( D => n1789, CK => n2054, Q => n_1024, QN 
                           => n1491);
   SWP_reg_2_inst : DFF_X1 port map( D => n1791, CK => n2047, Q => n1889, QN =>
                           n1493);
   SWP_reg_3_inst : DFF_X1 port map( D => n1790, CK => n2051, Q => n1934, QN =>
                           n1492);
   CANSAVE_reg_1_inst : DFF_X1 port map( D => n1796, CK => n2074, Q => n_1025, 
                           QN => n3284);
   CWP_reg_0_inst : DFF_X1 port map( D => n1788, CK => n2050, Q => CWP_0_port, 
                           QN => n1490);
   CWP_reg_1_inst : DFF_X1 port map( D => n1787, CK => n2051, Q => CWP_1_port, 
                           QN => n1489);
   CWP_reg_2_inst : DFF_X1 port map( D => n1786, CK => n2050, Q => CWP_2_port, 
                           QN => n1488);
   CWP_reg_3_inst : DFF_X1 port map( D => n1785, CK => n2050, Q => CWP_3_port, 
                           QN => n1487);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1656, CK => n2062, Q => 
                           n3118, QN => n1995);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1657, CK => n2062, Q => 
                           n3130, QN => n1994);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1658, CK => n2062, Q => 
                           n3142, QN => n1993);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1659, CK => n2062, Q => 
                           n3154, QN => n1992);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1660, CK => n2062, Q => 
                           n3166, QN => n1991);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1661, CK => n2062, Q => 
                           n3178, QN => n1990);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1662_port, CK => n2062, Q 
                           => n3190, QN => n1989);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1663_port, CK => n2062, Q 
                           => n3202, QN => n1988);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1664_port, CK => n2069, Q 
                           => n3111, QN => n1871);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1665_port, CK => n2069, Q 
                           => n3121, QN => n1917);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1666_port, CK => n2069, Q 
                           => n3133, QN => n1916);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1667, CK => n2069, Q => 
                           n3145, QN => n1915);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1668, CK => n2069, Q => 
                           n3157, QN => n1914);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1669, CK => n2069, Q => 
                           n3169, QN => n1913);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1670, CK => n2070, Q => 
                           n3181, QN => n1912);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1671, CK => n2070, Q => 
                           n3193, QN => n1911);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1672, CK => n2068, Q => 
                           n3069, QN => n1909);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1673, CK => n2068, Q => 
                           n3070, QN => n2012);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1674, CK => n2068, Q => 
                           n3071, QN => n2011);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1675, CK => n2068, Q => 
                           n3072, QN => n2010);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1676, CK => n2068, Q => 
                           n3073, QN => n2009);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1677, CK => n2068, Q => 
                           n3074, QN => n2008);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1678, CK => n2068, Q => 
                           n3075, QN => n2007);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1679, CK => n2068, Q => 
                           n3076, QN => n2006);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1680, CK => n2065, Q => 
                           n_1026, QN => n1839);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1681, CK => n2065, Q => 
                           n3231, QN => n1931);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1682, CK => n2065, Q => 
                           n3239, QN => n1930);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1683, CK => n2065, Q => 
                           n3247, QN => n1929);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1684, CK => n2065, Q => 
                           n3255, QN => n1928);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1685, CK => n2065, Q => 
                           n3263, QN => n1927);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1686, CK => n2065, Q => 
                           n3271, QN => n1926);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1687, CK => n2065, Q => 
                           n3279, QN => n1925);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1624, CK => n2064, Q => 
                           n3053, QN => n2027);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1625, CK => n2064, Q => 
                           n3054, QN => n2026);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1626, CK => n2064, Q => 
                           n3055, QN => n2025);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => n2064, Q => 
                           n3056, QN => n2024);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1628, CK => n2064, Q => 
                           n3057, QN => n2023);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1629, CK => n2064, Q => 
                           n3058, QN => n2022);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1630, CK => n2064, Q => 
                           n3059, QN => n2021);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1631, CK => n2065, Q => 
                           n3060, QN => n2020);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1632, CK => n2063, Q => 
                           n3110, QN => n1980);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1633, CK => n2063, Q => 
                           n3120, QN => n1979);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1634, CK => n2063, Q => 
                           n3132, QN => n1978);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1635, CK => n2063, Q => 
                           n3144, QN => n1977);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1636, CK => n2064, Q => 
                           n3156, QN => n1976);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1637, CK => n2064, Q => 
                           n3168, QN => n1975);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1638, CK => n2064, Q => 
                           n3180, QN => n1974);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1639, CK => n2064, Q => 
                           n3192, QN => n1973);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1640, CK => n2073, Q => 
                           n3061, QN => n1908);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1641, CK => n2073, Q => 
                           n3062, QN => n2019);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1642, CK => n2073, Q => 
                           n3063, QN => n2018);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1643, CK => n2073, Q => 
                           n3064, QN => n2017);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1644, CK => n2073, Q => 
                           n3065, QN => n2016);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1645, CK => n2073, Q => 
                           n3066, QN => n2015);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1646, CK => n2073, Q => 
                           n3067, QN => n2014);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1647, CK => n2073, Q => 
                           n3068, QN => n2013);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1648, CK => n2062, Q => 
                           n_1027, QN => n1815);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1649, CK => n2063, Q => 
                           n3229, QN => n1879);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1650, CK => n2063, Q => 
                           n3237, QN => n1878);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1651, CK => n2063, Q => 
                           n3245, QN => n1877);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1652, CK => n2063, Q => 
                           n3253, QN => n1876);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1653, CK => n2063, Q => 
                           n3261, QN => n1875);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1654, CK => n2063, Q => 
                           n3269, QN => n1874);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1655, CK => n2063, Q => 
                           n3277, QN => n1873);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1688, CK => n2051, Q => 
                           n3077, QN => n1996);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1689, CK => n2052, Q => 
                           n3078, QN => n1972);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1690, CK => n2052, Q => 
                           n3079, QN => n1971);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1691, CK => n2052, Q => 
                           n3080, QN => n1970);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1692, CK => n2052, Q => 
                           n3081, QN => n1969);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1693, CK => n2052, Q => 
                           n3082, QN => n1968);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1694, CK => n2052, Q => 
                           n3083, QN => n1967);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1695, CK => n2052, Q => 
                           n3084, QN => n1966);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1696, CK => n2052, Q => 
                           n3085, QN => n1872);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1697, CK => n2052, Q => 
                           n3086, QN => n1862);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1698, CK => n2052, Q => 
                           n3087, QN => n1860);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1699, CK => n2052, Q => 
                           n3088, QN => n1858);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1700, CK => n2053, Q => 
                           n3089, QN => n1856);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1701, CK => n2053, Q => 
                           n3090, QN => n1854);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1702, CK => n2053, Q => 
                           n3091, QN => n1852);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1703, CK => n2053, Q => 
                           n3092, QN => n1850);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1704, CK => n2073, Q => 
                           n3203, QN => n1848);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1705, CK => n2073, Q => 
                           n3205, QN => n1965);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1706, CK => n2074, Q => 
                           n3207, QN => n1963);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1707, CK => n2074, Q => 
                           n3209, QN => n1961);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1708, CK => n2074, Q => 
                           n3211, QN => n1959);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1709, CK => n2074, Q => 
                           n3213, QN => n1957);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1710, CK => n2074, Q => 
                           n3215, QN => n1955);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1711, CK => n2074, Q => 
                           n3217, QN => n1953);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1712, CK => n2053, Q => 
                           n_1028, QN => n1890);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1713, CK => n2053, Q => 
                           n_1029, QN => n1806);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1714, CK => n2053, Q => 
                           n_1030, QN => n1805);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1715, CK => n2053, Q => 
                           n_1031, QN => n1804);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1716, CK => n2053, Q => 
                           n_1032, QN => n1803);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1717, CK => n2053, Q => 
                           n_1033, QN => n1802);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1718, CK => n2053, Q => 
                           n_1034, QN => n1801);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1719, CK => n2054, Q => 
                           n_1035, QN => n1800);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1720, CK => n2054, Q => 
                           n3117, QN => n1880);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1721, CK => n2054, Q => 
                           n3129, QN => n1822);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1722, CK => n2054, Q => 
                           n3141, QN => n1821);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1723, CK => n2054, Q => 
                           n3153, QN => n1820);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1724, CK => n2054, Q => 
                           n3165, QN => n1819);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1725, CK => n2054, Q => 
                           n3177, QN => n1818);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1726, CK => n2054, Q => 
                           n3189, QN => n1817);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1727, CK => n2054, Q => 
                           n3201, QN => n1816);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1728, CK => n2068, Q => 
                           n3093, QN => n1932);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1729, CK => n2068, Q => 
                           n3094, QN => n1863);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1730, CK => n2068, Q => 
                           n3095, QN => n1861);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1731, CK => n2069, Q => 
                           n3096, QN => n1859);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1732, CK => n2069, Q => 
                           n3097, QN => n1857);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1733, CK => n2069, Q => 
                           n3098, QN => n1855);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1734, CK => n2069, Q => 
                           n3099, QN => n1853);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1735, CK => n2069, Q => 
                           n3100, QN => n1851);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1736, CK => n2065, Q => 
                           n3204, QN => n1849);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1737, CK => n2065, Q => 
                           n3206, QN => n1964);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1738, CK => n2066, Q => 
                           n3208, QN => n1962);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1739, CK => n2066, Q => 
                           n3210, QN => n1960);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1740, CK => n2066, Q => 
                           n3212, QN => n1958);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1741, CK => n2066, Q => 
                           n3214, QN => n1956);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1742, CK => n2066, Q => 
                           n3216, QN => n1954);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1743, CK => n2066, Q => 
                           n3218, QN => n1952);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1744, CK => n2051, Q => 
                           n3224, QN => n1910);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1745, CK => n2051, Q => 
                           n3232, QN => n1870);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1746, CK => n2051, Q => 
                           n3240, QN => n1869);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1747, CK => n2051, Q => 
                           n3248, QN => n1868);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1748, CK => n2051, Q => 
                           n3256, QN => n1867);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1749, CK => n2051, Q => 
                           n3264, QN => n1866);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1750, CK => n2051, Q => 
                           n3272, QN => n1865);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1751, CK => n2051, Q => 
                           n3280, QN => n1864);
   CWP_reg_4_inst : DFF_X1 port map( D => n1784, CK => n2050, Q => CWP_4_port, 
                           QN => n1486);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1496, CK => n2057, Q => 
                           n3116, QN => n1997);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1497, CK => n2057, Q => 
                           n3126, QN => n2004);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1498, CK => n2058, Q => 
                           n3138, QN => n2003);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1499, CK => n2058, Q => 
                           n3150, QN => n2002);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1500, CK => n2058, Q => 
                           n3162, QN => n2001);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1501, CK => n2058, Q => 
                           n3174, QN => n2000);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1502, CK => n2058, Q => 
                           n3186, QN => n1999);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1503, CK => n2058, Q => 
                           n3198, QN => n1998);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1504, CK => n2055, Q => 
                           n_1036, QN => n3113);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1505, CK => n2055, Q => 
                           n_1037, QN => n3123);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1506, CK => n2055, Q => 
                           n_1038, QN => n3135);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1507, CK => n2055, Q => 
                           n_1039, QN => n3147);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1508, CK => n2056, Q => 
                           n_1040, QN => n3159);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1509, CK => n2056, Q => 
                           n_1041, QN => n3171);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1510, CK => n2056, Q => 
                           n_1042, QN => n3183);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1511, CK => n2056, Q => 
                           n_1043, QN => n3195);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1512, CK => n2072, Q => 
                           n_1044, QN => n1807);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1513, CK => n2072, Q => 
                           n3127, QN => n1888);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1514, CK => n2072, Q => 
                           n3139, QN => n1887);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1515, CK => n2072, Q => 
                           n3151, QN => n1886);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1516, CK => n2072, Q => 
                           n3163, QN => n1885);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1517, CK => n2072, Q => 
                           n3175, QN => n1884);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1518, CK => n2072, Q => 
                           n3187, QN => n1883);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1519, CK => n2073, Q => 
                           n3199, QN => n1882);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1520, CK => n2056, Q => 
                           n_1045, QN => n3112);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1521, CK => n2056, Q => 
                           n_1046, QN => n3122);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1522, CK => n2056, Q => 
                           n_1047, QN => n3134);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1523, CK => n2056, Q => 
                           n_1048, QN => n3146);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1524, CK => n2056, Q => 
                           n_1049, QN => n3158);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1525, CK => n2056, Q => 
                           n_1050, QN => n3170);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1526, CK => n2056, Q => 
                           n_1051, QN => n3182);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1527, CK => n2057, Q => 
                           n_1052, QN => n3194);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n1528, CK => n2057, Q => 
                           n3115, QN => n1881);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n1529, CK => n2057, Q => 
                           n3125, QN => n1829);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n1530, CK => n2057, Q => 
                           n3137, QN => n1828);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n1531, CK => n2057, Q => 
                           n3149, QN => n1827);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n1532, CK => n2057, Q => 
                           n3161, QN => n1826);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n1533, CK => n2057, Q => 
                           n3173, QN => n1825);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n1534, CK => n2057, Q => 
                           n3185, QN => n1824);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n1535, CK => n2057, Q => 
                           n3197, QN => n1823);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1536, CK => n2070, Q => 
                           n_1053, QN => n3114);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1537, CK => n2070, Q => 
                           n_1054, QN => n3124);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1538, CK => n2070, Q => 
                           n_1055, QN => n3136);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1539, CK => n2070, Q => 
                           n_1056, QN => n3148);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1540, CK => n2070, Q => 
                           n_1057, QN => n3160);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1541, CK => n2070, Q => 
                           n_1058, QN => n3172);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1542, CK => n2070, Q => 
                           n_1059, QN => n3184);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1543, CK => n2070, Q => 
                           n_1060, QN => n3196);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1544, CK => n2066, Q => 
                           n3045, QN => n1907);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1545, CK => n2066, Q => 
                           n3046, QN => n2034);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1546, CK => n2066, Q => 
                           n3047, QN => n2033);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1547, CK => n2066, Q => 
                           n3048, QN => n2032);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1548, CK => n2066, Q => 
                           n3049, QN => n2031);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1549, CK => n2067, Q => 
                           n3050, QN => n2030);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1550, CK => n2067, Q => 
                           n3051, QN => n2029);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1551, CK => n2067, Q => 
                           n3052, QN => n2028);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1552, CK => n2054, Q => 
                           n3223, QN => n1901);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1553, CK => n2055, Q => 
                           n3230, QN => n1900);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1554, CK => n2055, Q => 
                           n3238, QN => n1899);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1555, CK => n2055, Q => 
                           n3246, QN => n1898);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1556, CK => n2055, Q => 
                           n3254, QN => n1897);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1557, CK => n2055, Q => 
                           n3262, QN => n1896);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1558, CK => n2055, Q => 
                           n3270, QN => n1895);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1559, CK => n2055, Q => 
                           n3278, QN => n1894);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1560, CK => n2061, Q => 
                           n1840, QN => n3221);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1561, CK => n2061, Q => 
                           n1841, QN => n3227);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1562, CK => n2061, Q => 
                           n1847, QN => n3235);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1563, CK => n2061, Q => 
                           n1846, QN => n3243);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1564, CK => n2061, Q => 
                           n1845, QN => n3251);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1565, CK => n2061, Q => 
                           n1844, QN => n3259);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1566, CK => n2062, Q => 
                           n1843, QN => n3267);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1567, CK => n2062, Q => 
                           n1842, QN => n3275);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1568, CK => n2060, Q => 
                           n_1061, QN => n1891);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1569, CK => n2060, Q => 
                           n_1062, QN => n1814);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1570, CK => n2060, Q => 
                           n_1063, QN => n1813);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1571, CK => n2060, Q => 
                           n_1064, QN => n1812);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1572, CK => n2060, Q => 
                           n_1065, QN => n1811);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1573, CK => n2060, Q => 
                           n_1066, QN => n1810);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1574, CK => n2060, Q => 
                           n_1067, QN => n1809);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1575, CK => n2060, Q => 
                           n_1068, QN => n1808);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1576, CK => n2071, Q => 
                           n2005, QN => n3222);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1577, CK => n2071, Q => 
                           n1893, QN => n3228);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1578, CK => n2071, Q => 
                           n1892, QN => n3236);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1579, CK => n2071, Q => 
                           n1906, QN => n3244);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1580, CK => n2072, Q => 
                           n1905, QN => n3252);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1581, CK => n2072, Q => 
                           n1904, QN => n3260);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1582, CK => n2072, Q => 
                           n1903, QN => n3268);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1583, CK => n2072, Q => 
                           n1902, QN => n3276);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1584, CK => n2060, Q => 
                           n_1069, QN => n1838);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1585, CK => n2060, Q => 
                           n_1070, QN => n1837);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1586, CK => n2060, Q => 
                           n_1071, QN => n1836);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1587, CK => n2061, Q => 
                           n_1072, QN => n1835);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1588, CK => n2061, Q => 
                           n_1073, QN => n1834);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1589, CK => n2061, Q => 
                           n_1074, QN => n1833);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1590, CK => n2061, Q => 
                           n_1075, QN => n1832);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1591, CK => n2061, Q => 
                           n_1076, QN => n1831);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1592, CK => n2059, Q => 
                           n1935, QN => n3220);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1593, CK => n2059, Q => 
                           n1937, QN => n3226);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1594, CK => n2059, Q => 
                           n1943, QN => n3234);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1595, CK => n2059, Q => 
                           n1942, QN => n3242);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1596, CK => n2059, Q => 
                           n1941, QN => n3250);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1597, CK => n2059, Q => 
                           n1940, QN => n3258);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1598, CK => n2059, Q => 
                           n1939, QN => n3266);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1599, CK => n2059, Q => 
                           n1938, QN => n3274);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1600, CK => n2070, Q => 
                           n_1077, QN => n3036);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1601, CK => n2071, Q => 
                           n_1078, QN => n3035);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1602, CK => n2071, Q => 
                           n_1079, QN => n3034);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1603, CK => n2071, Q => 
                           n_1080, QN => n3033);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1604, CK => n2071, Q => 
                           n_1081, QN => n3032);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1605, CK => n2071, Q => 
                           n_1082, QN => n3031);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1606, CK => n2071, Q => 
                           n_1083, QN => n3030);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1607, CK => n2071, Q => 
                           n_1084, QN => n3029);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1608, CK => n2067, Q => 
                           n_1085, QN => n1799);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1609, CK => n2067, Q => 
                           n3128, QN => n1987);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1610, CK => n2067, Q => 
                           n3140, QN => n1986);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1611, CK => n2067, Q => 
                           n3152, QN => n1985);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1612, CK => n2067, Q => 
                           n3164, QN => n1984);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1613, CK => n2067, Q => 
                           n3176, QN => n1983);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1614, CK => n2067, Q => 
                           n3188, QN => n1982);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1615, CK => n2067, Q => 
                           n3200, QN => n1981);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1616, CK => n2058, Q => 
                           n_1086, QN => n3109);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1617, CK => n2058, Q => 
                           n_1087, QN => n3119);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1618, CK => n2058, Q => 
                           n_1088, QN => n3131);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1619, CK => n2058, Q => 
                           n_1089, QN => n3143);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1620, CK => n2058, Q => 
                           n_1090, QN => n3155);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1621, CK => n2059, Q => 
                           n_1091, QN => n3167);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1622, CK => n2059, Q => 
                           n_1092, QN => n3179);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1623, CK => n2059, Q => 
                           n_1093, QN => n3191);
   r121 : WINDOWED_REGISTER_FILE_DW01_addsub_0_DW01_addsub_2 port map( A(4) => 
                           CWP_4_port, A(3) => CWP_3_port, A(2) => CWP_2_port, 
                           A(1) => CWP_1_port, A(0) => CWP_0_port, B(4) => n10,
                           B(3) => U3_U22_Z_3, B(2) => U3_U22_Z_2, B(1) => 
                           U3_U22_Z_1, B(0) => U3_U22_Z_0, CI => n10, ADD_SUB 
                           => U3_U23_Z_0, SUM(4) => N1666, SUM(3) => N1665, 
                           SUM(2) => N1664, SUM(1) => N1663, SUM(0) => N1662, 
                           CO => n_1094);
   OUT2_tri_0_inst : TBUF_X1 port map( A => n1264, EN => n1257, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n1263, EN => n1257, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n1262, EN => n1257, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n1261, EN => n1257, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n1260, EN => n1257, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n1259, EN => n1257, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n1258, EN => n1257, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n1256, EN => n1257, Z => OUT2(7));
   OUT1_tri_0_inst : TBUF_X1 port map( A => n1255, EN => n1248, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n1254, EN => n1248, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n1253, EN => n1248, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n1252, EN => n1248, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n1251, EN => n1248, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n1250, EN => n1248, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n1249, EN => n1248, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n1247, EN => n1248, Z => OUT1(7));
   TO_MEM_tri_0_inst : TBUF_X1 port map( A => n1273, EN => n1266, Z => 
                           TO_MEM(0));
   TO_MEM_tri_1_inst : TBUF_X1 port map( A => n1272, EN => n1266, Z => 
                           TO_MEM(1));
   TO_MEM_tri_2_inst : TBUF_X1 port map( A => n1271, EN => n1266, Z => 
                           TO_MEM(2));
   TO_MEM_tri_3_inst : TBUF_X1 port map( A => n1270, EN => n1266, Z => 
                           TO_MEM(3));
   TO_MEM_tri_4_inst : TBUF_X1 port map( A => n1269, EN => n1266, Z => 
                           TO_MEM(4));
   TO_MEM_tri_5_inst : TBUF_X1 port map( A => n1268, EN => n1266, Z => 
                           TO_MEM(5));
   TO_MEM_tri_6_inst : TBUF_X1 port map( A => n1267, EN => n1266, Z => 
                           TO_MEM(6));
   TO_MEM_tri_7_inst : TBUF_X1 port map( A => n1265, EN => n1266, Z => 
                           TO_MEM(7));
   U1477 : AOI221_X1 port map( B1 => n2562, B2 => n3062, C1 => n2563, C2 => 
                           n3229, A => n2725, ZN => n2722);
   U1478 : AOI221_X1 port map( B1 => n2557, B2 => n1893, C1 => n2558, C2 => 
                           n3127, A => n2724, ZN => n2723);
   U1479 : AOI221_X1 port map( B1 => n2562, B2 => n3070, C1 => n2563, C2 => 
                           n3231, A => n2721, ZN => n2718);
   U1480 : AOI221_X1 port map( B1 => n2557, B2 => n3128, C1 => n2558, C2 => 
                           n3046, A => n2720, ZN => n2719);
   U1481 : AOI221_X1 port map( B1 => n2562, B2 => n3130, C1 => n2563, C2 => 
                           n3121, A => n2717, ZN => n2713);
   U1482 : AOI221_X1 port map( B1 => n2557, B2 => n1937, C1 => n2558, C2 => 
                           n3125, A => n2716, ZN => n2714);
   U1483 : AOI221_X1 port map( B1 => n2562, B2 => n3054, C1 => n2563, C2 => 
                           n3120, A => n2712, ZN => n2708);
   U1484 : AOI221_X1 port map( B1 => n2557, B2 => n1841, C1 => n2558, C2 => 
                           n3126, A => n2711, ZN => n2709);
   U1485 : AOI221_X1 port map( B1 => n2562, B2 => n3063, C1 => n2563, C2 => 
                           n3237, A => n2700, ZN => n2697);
   U1486 : AOI221_X1 port map( B1 => n2557, B2 => n1892, C1 => n2558, C2 => 
                           n3139, A => n2699, ZN => n2698);
   U1487 : AOI221_X1 port map( B1 => n2562, B2 => n3071, C1 => n2563, C2 => 
                           n3239, A => n2696, ZN => n2693);
   U1488 : AOI221_X1 port map( B1 => n2557, B2 => n3140, C1 => n2558, C2 => 
                           n3047, A => n2695, ZN => n2694);
   U1489 : AOI221_X1 port map( B1 => n2818, B2 => n1945, C1 => n2819, C2 => 
                           n3102, A => n2962, ZN => n2938);
   U1490 : AOI221_X1 port map( B1 => n2818, B2 => n1946, C1 => n2819, C2 => 
                           n3103, A => n2937, ZN => n2915);
   U1491 : AOI221_X1 port map( B1 => n2582, B2 => n1945, C1 => n2583, C2 => 
                           n3102, A => n2726, ZN => n2702);
   U1492 : AOI221_X1 port map( B1 => n2582, B2 => n1946, C1 => n2583, C2 => 
                           n3103, A => n2701, ZN => n2679);
   U1493 : AOI221_X1 port map( B1 => n2582, B2 => n1947, C1 => n2583, C2 => 
                           n3107, A => n2609, ZN => n2587);
   U1494 : AOI221_X1 port map( B1 => n2582, B2 => n1948, C1 => n2583, C2 => 
                           n3106, A => n2632, ZN => n2610);
   U1495 : AOI221_X1 port map( B1 => n2582, B2 => n1949, C1 => n2583, C2 => 
                           n3105, A => n2655, ZN => n2633);
   U1496 : AOI221_X1 port map( B1 => n2582, B2 => n1950, C1 => n2583, C2 => 
                           n3104, A => n2678, ZN => n2656);
   U1497 : NOR3_X2 port map( A1 => n2755, A2 => n2753, A3 => n2738, ZN => n2582
                           );
   U1498 : AOI221_X1 port map( B1 => n2818, B2 => n1947, C1 => n2819, C2 => 
                           n3107, A => n2845, ZN => n2823);
   U1499 : AOI221_X1 port map( B1 => n2818, B2 => n1948, C1 => n2819, C2 => 
                           n3106, A => n2868, ZN => n2846);
   U1500 : AOI221_X1 port map( B1 => n2818, B2 => n1949, C1 => n2819, C2 => 
                           n3105, A => n2891, ZN => n2869);
   U1501 : AOI221_X1 port map( B1 => n2818, B2 => n1950, C1 => n2819, C2 => 
                           n3104, A => n2914, ZN => n2892);
   U1502 : NOR3_X2 port map( A1 => n2990, A2 => n2988, A3 => n2973, ZN => n2818
                           );
   U1503 : NOR3_X2 port map( A1 => n2753, A2 => ADD_RD2(1), A3 => n2738, ZN => 
                           n2583);
   U1504 : NOR3_X2 port map( A1 => n2988, A2 => ADD_RD1(1), A3 => n2973, ZN => 
                           n2819);
   U1505 : NAND2_X2 port map( A1 => FROM_MEM(6), A2 => n2405, ZN => n2191);
   U1506 : NAND3_X2 port map( A1 => n3006, A2 => n3005, A3 => n3004, ZN => 
                           n2801);
   U1507 : NAND2_X2 port map( A1 => FROM_MEM(5), A2 => n2405, ZN => n2190);
   U1508 : NAND3_X2 port map( A1 => n3002, A2 => n3003, A3 => n3004, ZN => 
                           n2796);
   U1509 : NAND2_X2 port map( A1 => FROM_MEM(4), A2 => n2405, ZN => n2189);
   U1510 : NAND3_X2 port map( A1 => n3003, A2 => n3006, A3 => n3004, ZN => 
                           n2802);
   U1511 : NAND2_X2 port map( A1 => FROM_MEM(3), A2 => n2405, ZN => n2188);
   U1512 : NAND3_X2 port map( A1 => n3002, A2 => n3005, A3 => n3004, ZN => 
                           n2797);
   U1513 : INV_X2 port map( A => n2747, ZN => n2557);
   U1514 : NAND2_X2 port map( A1 => FROM_MEM(2), A2 => n2405, ZN => n2187);
   U1515 : INV_X1 port map( A => n2982, ZN => n2043);
   U1516 : INV_X2 port map( A => n2745, ZN => n2562);
   U1517 : NAND2_X2 port map( A1 => FROM_MEM(1), A2 => n2405, ZN => n2186);
   U1518 : NAND3_X2 port map( A1 => n2768, A2 => n2771, A3 => n2770, ZN => 
                           n2565);
   U1519 : NAND3_X2 port map( A1 => n2772, A2 => n2767, A3 => n2769, ZN => 
                           n2560);
   U1520 : INV_X1 port map( A => n2980, ZN => n2044);
   U1521 : NAND3_X2 port map( A1 => n1889, A2 => n1830, A3 => n1495, ZN => 
                           n2274);
   U1522 : INV_X2 port map( A => n2746, ZN => n2558);
   U1523 : NAND2_X2 port map( A1 => FROM_MEM(0), A2 => n2405, ZN => n2185);
   U1524 : NAND3_X2 port map( A1 => n2768, A2 => n2771, A3 => n2769, ZN => 
                           n2566);
   U1525 : INV_X1 port map( A => n2981, ZN => n2045);
   U1526 : INV_X2 port map( A => n2744, ZN => n2563);
   U1527 : NAND2_X2 port map( A1 => FROM_MEM(7), A2 => n2405, ZN => n2192);
   U1528 : NAND3_X2 port map( A1 => n2772, A2 => n2771, A3 => n2769, ZN => 
                           n2561);
   U1529 : AOI21_X4 port map( B1 => n2139, B2 => n2409, A => RESET, ZN => n2181
                           );
   U1530 : INV_X1 port map( A => n2979, ZN => n2046);
   U1531 : BUF_X1 port map( A => CLK, Z => n2090);
   U1532 : BUF_X1 port map( A => CLK, Z => n2089);
   U1533 : BUF_X1 port map( A => n2082, Z => n2059);
   U1534 : BUF_X1 port map( A => n2076, Z => n2071);
   U1535 : BUF_X1 port map( A => n2082, Z => n2060);
   U1536 : BUF_X1 port map( A => n2081, Z => n2061);
   U1537 : BUF_X1 port map( A => n2078, Z => n2067);
   U1538 : BUF_X1 port map( A => n2076, Z => n2072);
   U1539 : BUF_X1 port map( A => n2084, Z => n2056);
   U1540 : BUF_X1 port map( A => n2084, Z => n2055);
   U1541 : BUF_X1 port map( A => n2083, Z => n2058);
   U1542 : BUF_X1 port map( A => n2083, Z => n2057);
   U1543 : BUF_X1 port map( A => n2079, Z => n2066);
   U1544 : BUF_X1 port map( A => n2085, Z => n2053);
   U1545 : BUF_X1 port map( A => n2086, Z => n2052);
   U1546 : BUF_X1 port map( A => n2075, Z => n2073);
   U1547 : BUF_X1 port map( A => n2080, Z => n2063);
   U1548 : BUF_X1 port map( A => n2080, Z => n2064);
   U1549 : BUF_X1 port map( A => n2079, Z => n2065);
   U1550 : BUF_X1 port map( A => n2078, Z => n2068);
   U1551 : BUF_X1 port map( A => n2077, Z => n2070);
   U1552 : BUF_X1 port map( A => n2077, Z => n2069);
   U1553 : BUF_X1 port map( A => n2081, Z => n2062);
   U1554 : BUF_X1 port map( A => n2086, Z => n2051);
   U1555 : BUF_X1 port map( A => n2085, Z => n2054);
   U1556 : BUF_X1 port map( A => n2087, Z => n2049);
   U1557 : BUF_X1 port map( A => n2088, Z => n2048);
   U1558 : BUF_X1 port map( A => n2087, Z => n2050);
   U1559 : BUF_X1 port map( A => n2088, Z => n2047);
   U1560 : BUF_X1 port map( A => n2075, Z => n2074);
   U1561 : BUF_X1 port map( A => n2090, Z => n2082);
   U1562 : BUF_X1 port map( A => n2089, Z => n2084);
   U1563 : BUF_X1 port map( A => n2090, Z => n2083);
   U1564 : BUF_X1 port map( A => n2090, Z => n2080);
   U1565 : BUF_X1 port map( A => n2090, Z => n2079);
   U1566 : BUF_X1 port map( A => n2090, Z => n2081);
   U1567 : BUF_X1 port map( A => n2089, Z => n2086);
   U1568 : BUF_X1 port map( A => n2089, Z => n2085);
   U1569 : BUF_X1 port map( A => n2089, Z => n2087);
   U1570 : BUF_X1 port map( A => n2089, Z => n2088);
   U1571 : BUF_X1 port map( A => n2091, Z => n2076);
   U1572 : BUF_X1 port map( A => n2091, Z => n2078);
   U1573 : BUF_X1 port map( A => n2091, Z => n2077);
   U1574 : BUF_X1 port map( A => n2091, Z => n2075);
   U1575 : BUF_X1 port map( A => CLK, Z => n2091);
   U1576 : NAND2_X1 port map( A1 => n2092, A2 => n2093, ZN => n1797);
   U1577 : XOR2_X1 port map( A => n2094, B => n3285, Z => n2092);
   U1578 : NAND3_X1 port map( A1 => n2095, A2 => n2093, A3 => n2096, ZN => 
                           n1796);
   U1579 : XNOR2_X1 port map( A => n3284, B => n2097, ZN => n2096);
   U1580 : OAI21_X1 port map( B1 => CALL, B2 => n3285, A => n2098, ZN => n2097)
                           ;
   U1581 : NAND3_X1 port map( A1 => CALL, A2 => n3285, A3 => n2098, ZN => n2095
                           );
   U1582 : INV_X1 port map( A => n2094, ZN => n2098);
   U1583 : NAND2_X1 port map( A1 => n2099, A2 => n2093, ZN => n1795);
   U1584 : XOR2_X1 port map( A => n2094, B => n3281, Z => n2099);
   U1585 : NAND2_X1 port map( A1 => n2100, A2 => n2093, ZN => n1794);
   U1586 : XNOR2_X1 port map( A => n3282, B => n2101, ZN => n2100);
   U1587 : NOR2_X1 port map( A1 => n2102, A2 => n2094, ZN => n2101);
   U1588 : XNOR2_X1 port map( A => n3281, B => n2103, ZN => n2102);
   U1589 : MUX2_X1 port map( A => n2104, B => n2105, S => n1495, Z => n1793);
   U1590 : NAND2_X1 port map( A1 => n2106, A2 => n2107, ZN => n2105);
   U1591 : INV_X1 port map( A => n2108, ZN => n2104);
   U1592 : OAI222_X1 port map( A1 => n1494, A2 => n2109, B1 => n1495, B2 => 
                           n2110, C1 => n2111, C2 => n2106, ZN => n1792);
   U1593 : MUX2_X1 port map( A => n2106, B => n2107, S => n1494, Z => n2110);
   U1594 : INV_X1 port map( A => n2112, ZN => n2109);
   U1595 : OAI222_X1 port map( A1 => n2107, A2 => n2113, B1 => n1493, B2 => 
                           n2114, C1 => n2106, C2 => n2115, ZN => n1791);
   U1596 : AOI221_X1 port map( B1 => n2116, B2 => n1494, C1 => n2117, C2 => 
                           n2111, A => n2112, ZN => n2114);
   U1597 : OAI21_X1 port map( B1 => n1798, B2 => n2107, A => n2108, ZN => n2112
                           );
   U1598 : MUX2_X1 port map( A => n2118, B => n2119, S => n1492, Z => n1790);
   U1599 : OAI22_X1 port map( A1 => n2106, A2 => n2115, B1 => n2107, B2 => 
                           n2120, ZN => n2119);
   U1600 : OAI211_X1 port map( C1 => n1491, C2 => n2121, A => n2122, B => n2123
                           , ZN => n1789);
   U1601 : OAI21_X1 port map( B1 => n2124, B2 => n2125, A => n2116, ZN => n2123
                           );
   U1602 : INV_X1 port map( A => n2107, ZN => n2116);
   U1603 : INV_X1 port map( A => n2126, ZN => n2124);
   U1604 : OAI21_X1 port map( B1 => n2127, B2 => n2128, A => n2117, ZN => n2122
                           );
   U1605 : INV_X1 port map( A => n2106, ZN => n2117);
   U1606 : INV_X1 port map( A => n2118, ZN => n2121);
   U1607 : OAI221_X1 port map( B1 => n2129, B2 => n2107, C1 => n2130, C2 => 
                           n2106, A => n2108, ZN => n2118);
   U1608 : NAND2_X1 port map( A1 => n2131, A2 => n2108, ZN => n2106);
   U1609 : OAI21_X1 port map( B1 => CALL, B2 => n2132, A => n2133, ZN => n2131)
                           ;
   U1610 : NAND2_X1 port map( A1 => n2134, A2 => n2108, ZN => n2107);
   U1611 : NAND3_X1 port map( A1 => n2135, A2 => n2093, A3 => n2136, ZN => 
                           n2108);
   U1612 : NAND3_X1 port map( A1 => n2137, A2 => n2115, A3 => n2138, ZN => 
                           n2136);
   U1613 : NAND4_X1 port map( A1 => ENABLE, A2 => n2139, A3 => n2140, A4 => 
                           n2141, ZN => n2135);
   U1614 : OAI21_X1 port map( B1 => n2142, B2 => n2143, A => n2144, ZN => n2140
                           );
   U1615 : OAI22_X1 port map( A1 => RESET, A2 => n1266, B1 => n2144, B2 => 
                           n2132, ZN => n2134);
   U1616 : OAI22_X1 port map( A1 => n1490, A2 => n2145, B1 => n2146, B2 => 
                           n2147, ZN => n1788);
   U1617 : OAI22_X1 port map( A1 => n1489, A2 => n2145, B1 => n2146, B2 => 
                           n2148, ZN => n1787);
   U1618 : OAI22_X1 port map( A1 => n1488, A2 => n2145, B1 => n2146, B2 => 
                           n2149, ZN => n1786);
   U1619 : OAI22_X1 port map( A1 => n1487, A2 => n2145, B1 => n2146, B2 => 
                           n2150, ZN => n1785);
   U1620 : OAI22_X1 port map( A1 => n1486, A2 => n2145, B1 => n2146, B2 => 
                           n2151, ZN => n1784);
   U1621 : NAND2_X1 port map( A1 => n2093, A2 => n2145, ZN => n2146);
   U1622 : OAI211_X1 port map( C1 => n2115, C2 => n2152, A => n2094, B => n2093
                           , ZN => n2145);
   U1623 : NAND3_X1 port map( A1 => ENABLE, A2 => n2139, A3 => n2153, ZN => 
                           n2094);
   U1624 : MUX2_X1 port map( A => n2154, B => n2155, S => CALL, Z => n2153);
   U1625 : NAND2_X1 port map( A1 => n2138, A2 => n2137, ZN => n2152);
   U1626 : OAI22_X1 port map( A1 => n3273, A2 => n2156, B1 => n2157, B2 => 
                           n2158, ZN => n1783);
   U1627 : OAI22_X1 port map( A1 => n3265, A2 => n2156, B1 => n2157, B2 => 
                           n2159, ZN => n1782);
   U1628 : OAI22_X1 port map( A1 => n3257, A2 => n2156, B1 => n2157, B2 => 
                           n2160, ZN => n1781);
   U1629 : OAI22_X1 port map( A1 => n3249, A2 => n2156, B1 => n2157, B2 => 
                           n2161, ZN => n1780);
   U1630 : OAI22_X1 port map( A1 => n3241, A2 => n2156, B1 => n2157, B2 => 
                           n2162, ZN => n1779);
   U1631 : OAI22_X1 port map( A1 => n3233, A2 => n2156, B1 => n2157, B2 => 
                           n2163, ZN => n1778);
   U1632 : OAI22_X1 port map( A1 => n3225, A2 => n2156, B1 => n2157, B2 => 
                           n2164, ZN => n1777);
   U1633 : OAI22_X1 port map( A1 => n3219, A2 => n2156, B1 => n2157, B2 => 
                           n2165, ZN => n1776);
   U1634 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2166, A3 => ADD_WR(1), ZN
                           => n2157);
   U1635 : NAND2_X1 port map( A1 => n2093, A2 => n2167, ZN => n2156);
   U1636 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2168, A3 => ADD_WR(1), ZN
                           => n2167);
   U1637 : OAI22_X1 port map( A1 => n3037, A2 => n2169, B1 => n2158, B2 => 
                           n2170, ZN => n1775);
   U1638 : OAI22_X1 port map( A1 => n3038, A2 => n2169, B1 => n2159, B2 => 
                           n2170, ZN => n1774);
   U1639 : OAI22_X1 port map( A1 => n3039, A2 => n2169, B1 => n2160, B2 => 
                           n2170, ZN => n1773);
   U1640 : OAI22_X1 port map( A1 => n3040, A2 => n2169, B1 => n2161, B2 => 
                           n2170, ZN => n1772);
   U1641 : OAI22_X1 port map( A1 => n3041, A2 => n2169, B1 => n2162, B2 => 
                           n2170, ZN => n1771);
   U1642 : OAI22_X1 port map( A1 => n3042, A2 => n2169, B1 => n2163, B2 => 
                           n2170, ZN => n1770);
   U1643 : OAI22_X1 port map( A1 => n3043, A2 => n2169, B1 => n2164, B2 => 
                           n2170, ZN => n1769);
   U1644 : OAI22_X1 port map( A1 => n3044, A2 => n2169, B1 => n2165, B2 => 
                           n2170, ZN => n1768);
   U1645 : NAND3_X1 port map( A1 => n2166, A2 => n2171, A3 => ADD_WR(1), ZN => 
                           n2170);
   U1646 : NAND2_X1 port map( A1 => n2093, A2 => n2172, ZN => n2169);
   U1647 : NAND3_X1 port map( A1 => n2168, A2 => n2171, A3 => ADD_WR(1), ZN => 
                           n2172);
   U1648 : OAI22_X1 port map( A1 => n2173, A2 => n2036, B1 => n2158, B2 => 
                           n2174, ZN => n1767);
   U1649 : OAI22_X1 port map( A1 => n2173, A2 => n2037, B1 => n2159, B2 => 
                           n2174, ZN => n1766);
   U1650 : OAI22_X1 port map( A1 => n2173, A2 => n2038, B1 => n2160, B2 => 
                           n2174, ZN => n1765);
   U1651 : OAI22_X1 port map( A1 => n2173, A2 => n2039, B1 => n2161, B2 => 
                           n2174, ZN => n1764);
   U1652 : OAI22_X1 port map( A1 => n2173, A2 => n2040, B1 => n2162, B2 => 
                           n2174, ZN => n1763);
   U1653 : OAI22_X1 port map( A1 => n2173, A2 => n2041, B1 => n2163, B2 => 
                           n2174, ZN => n1762);
   U1654 : OAI22_X1 port map( A1 => n2173, A2 => n2042, B1 => n2164, B2 => 
                           n2174, ZN => n1761);
   U1655 : OAI22_X1 port map( A1 => n2173, A2 => n2035, B1 => n2165, B2 => 
                           n2174, ZN => n1760);
   U1656 : NAND3_X1 port map( A1 => n2166, A2 => n2175, A3 => ADD_WR(0), ZN => 
                           n2174);
   U1657 : NAND2_X1 port map( A1 => n2093, A2 => n2176, ZN => n2173);
   U1658 : NAND3_X1 port map( A1 => n2168, A2 => n2175, A3 => ADD_WR(0), ZN => 
                           n2176);
   U1659 : OAI22_X1 port map( A1 => n2177, A2 => n1918, B1 => n2158, B2 => 
                           n2178, ZN => n1759);
   U1660 : OAI22_X1 port map( A1 => n2177, A2 => n1919, B1 => n2159, B2 => 
                           n2178, ZN => n1758);
   U1661 : OAI22_X1 port map( A1 => n2177, A2 => n1920, B1 => n2160, B2 => 
                           n2178, ZN => n1757);
   U1662 : OAI22_X1 port map( A1 => n2177, A2 => n1921, B1 => n2161, B2 => 
                           n2178, ZN => n1756);
   U1663 : OAI22_X1 port map( A1 => n2177, A2 => n1922, B1 => n2162, B2 => 
                           n2178, ZN => n1755);
   U1664 : OAI22_X1 port map( A1 => n2177, A2 => n1923, B1 => n2163, B2 => 
                           n2178, ZN => n1754);
   U1665 : OAI22_X1 port map( A1 => n2177, A2 => n1924, B1 => n2164, B2 => 
                           n2178, ZN => n1753);
   U1666 : OAI22_X1 port map( A1 => n2177, A2 => n1933, B1 => n2165, B2 => 
                           n2178, ZN => n1752);
   U1667 : NAND3_X1 port map( A1 => n2171, A2 => n2175, A3 => n2166, ZN => 
                           n2178);
   U1668 : AND2_X1 port map( A1 => n2168, A2 => n2093, ZN => n2166);
   U1669 : NAND2_X1 port map( A1 => n2093, A2 => n2179, ZN => n2177);
   U1670 : NAND3_X1 port map( A1 => n2171, A2 => n2175, A3 => n2168, ZN => 
                           n2179);
   U1671 : NOR2_X1 port map( A1 => n2180, A2 => n2181, ZN => n2168);
   U1672 : OAI222_X1 port map( A1 => n2182, A2 => n1864, B1 => n2158, B2 => 
                           n2183, C1 => n2184, C2 => n2185, ZN => n1751);
   U1673 : OAI222_X1 port map( A1 => n2182, A2 => n1865, B1 => n2159, B2 => 
                           n2183, C1 => n2184, C2 => n2186, ZN => n1750);
   U1674 : OAI222_X1 port map( A1 => n2182, A2 => n1866, B1 => n2160, B2 => 
                           n2183, C1 => n2184, C2 => n2187, ZN => n1749);
   U1675 : OAI222_X1 port map( A1 => n2182, A2 => n1867, B1 => n2161, B2 => 
                           n2183, C1 => n2184, C2 => n2188, ZN => n1748);
   U1676 : OAI222_X1 port map( A1 => n2182, A2 => n1868, B1 => n2162, B2 => 
                           n2183, C1 => n2184, C2 => n2189, ZN => n1747);
   U1677 : OAI222_X1 port map( A1 => n2182, A2 => n1869, B1 => n2163, B2 => 
                           n2183, C1 => n2184, C2 => n2190, ZN => n1746);
   U1678 : OAI222_X1 port map( A1 => n2182, A2 => n1870, B1 => n2164, B2 => 
                           n2183, C1 => n2184, C2 => n2191, ZN => n1745);
   U1679 : OAI222_X1 port map( A1 => n2182, A2 => n1910, B1 => n2165, B2 => 
                           n2183, C1 => n2184, C2 => n2192, ZN => n1744);
   U1680 : NAND3_X1 port map( A1 => n2193, A2 => n2194, A3 => n2195, ZN => 
                           n2183);
   U1681 : AND2_X1 port map( A1 => n2193, A2 => n2196, ZN => n2182);
   U1682 : OAI21_X1 port map( B1 => n2197, B2 => n2198, A => n2199, ZN => n2196
                           );
   U1683 : INV_X1 port map( A => n2184, ZN => n2193);
   U1684 : OAI21_X1 port map( B1 => n2200, B2 => n2201, A => n2202, ZN => n2184
                           );
   U1685 : OAI222_X1 port map( A1 => n2158, A2 => n2203, B1 => n2204, B2 => 
                           n1952, C1 => n2185, C2 => n2205, ZN => n1743);
   U1686 : OAI222_X1 port map( A1 => n2159, A2 => n2203, B1 => n2204, B2 => 
                           n1954, C1 => n2186, C2 => n2205, ZN => n1742);
   U1687 : OAI222_X1 port map( A1 => n2160, A2 => n2203, B1 => n2204, B2 => 
                           n1956, C1 => n2187, C2 => n2205, ZN => n1741);
   U1688 : OAI222_X1 port map( A1 => n2161, A2 => n2203, B1 => n2204, B2 => 
                           n1958, C1 => n2188, C2 => n2205, ZN => n1740);
   U1689 : OAI222_X1 port map( A1 => n2162, A2 => n2203, B1 => n2204, B2 => 
                           n1960, C1 => n2189, C2 => n2205, ZN => n1739);
   U1690 : OAI222_X1 port map( A1 => n2163, A2 => n2203, B1 => n2204, B2 => 
                           n1962, C1 => n2190, C2 => n2205, ZN => n1738);
   U1691 : OAI222_X1 port map( A1 => n2164, A2 => n2203, B1 => n2204, B2 => 
                           n1964, C1 => n2191, C2 => n2205, ZN => n1737);
   U1692 : OAI222_X1 port map( A1 => n2165, A2 => n2203, B1 => n2204, B2 => 
                           n1849, C1 => n2192, C2 => n2205, ZN => n1736);
   U1693 : AND2_X1 port map( A1 => n2206, A2 => n2207, ZN => n2204);
   U1694 : OAI21_X1 port map( B1 => n2198, B2 => n2208, A => n2199, ZN => n2207
                           );
   U1695 : NAND3_X1 port map( A1 => n2209, A2 => n2195, A3 => n2206, ZN => 
                           n2203);
   U1696 : INV_X1 port map( A => n2205, ZN => n2206);
   U1697 : OAI21_X1 port map( B1 => n2210, B2 => n2201, A => n2202, ZN => n2205
                           );
   U1698 : OAI222_X1 port map( A1 => n2158, A2 => n2211, B1 => n2212, B2 => 
                           n1851, C1 => n2213, C2 => n2185, ZN => n1735);
   U1699 : OAI222_X1 port map( A1 => n2159, A2 => n2211, B1 => n2212, B2 => 
                           n1853, C1 => n2213, C2 => n2186, ZN => n1734);
   U1700 : OAI222_X1 port map( A1 => n2160, A2 => n2211, B1 => n2212, B2 => 
                           n1855, C1 => n2213, C2 => n2187, ZN => n1733);
   U1701 : OAI222_X1 port map( A1 => n2161, A2 => n2211, B1 => n2212, B2 => 
                           n1857, C1 => n2213, C2 => n2188, ZN => n1732);
   U1702 : OAI222_X1 port map( A1 => n2162, A2 => n2211, B1 => n2212, B2 => 
                           n1859, C1 => n2213, C2 => n2189, ZN => n1731);
   U1703 : OAI222_X1 port map( A1 => n2163, A2 => n2211, B1 => n2212, B2 => 
                           n1861, C1 => n2213, C2 => n2190, ZN => n1730);
   U1704 : OAI222_X1 port map( A1 => n2164, A2 => n2211, B1 => n2212, B2 => 
                           n1863, C1 => n2213, C2 => n2191, ZN => n1729);
   U1705 : OAI222_X1 port map( A1 => n2165, A2 => n2211, B1 => n2212, B2 => 
                           n1932, C1 => n2213, C2 => n2192, ZN => n1728);
   U1706 : INV_X1 port map( A => n2214, ZN => n2213);
   U1707 : AND2_X1 port map( A1 => n2215, A2 => n2214, ZN => n2212);
   U1708 : OAI21_X1 port map( B1 => n2198, B2 => n2216, A => n2199, ZN => n2215
                           );
   U1709 : NAND3_X1 port map( A1 => n2195, A2 => n2214, A3 => n2217, ZN => 
                           n2211);
   U1710 : OAI21_X1 port map( B1 => n2218, B2 => n2219, A => n2181, ZN => n2214
                           );
   U1711 : OAI222_X1 port map( A1 => n2158, A2 => n2220, B1 => n2221, B2 => 
                           n1816, C1 => n2222, C2 => n2185, ZN => n1727);
   U1712 : OAI222_X1 port map( A1 => n2159, A2 => n2220, B1 => n2221, B2 => 
                           n1817, C1 => n2222, C2 => n2186, ZN => n1726);
   U1713 : OAI222_X1 port map( A1 => n2160, A2 => n2220, B1 => n2221, B2 => 
                           n1818, C1 => n2222, C2 => n2187, ZN => n1725);
   U1714 : OAI222_X1 port map( A1 => n2161, A2 => n2220, B1 => n2221, B2 => 
                           n1819, C1 => n2222, C2 => n2188, ZN => n1724);
   U1715 : OAI222_X1 port map( A1 => n2162, A2 => n2220, B1 => n2221, B2 => 
                           n1820, C1 => n2222, C2 => n2189, ZN => n1723);
   U1716 : OAI222_X1 port map( A1 => n2163, A2 => n2220, B1 => n2221, B2 => 
                           n1821, C1 => n2222, C2 => n2190, ZN => n1722);
   U1717 : OAI222_X1 port map( A1 => n2164, A2 => n2220, B1 => n2221, B2 => 
                           n1822, C1 => n2222, C2 => n2191, ZN => n1721);
   U1718 : OAI222_X1 port map( A1 => n2165, A2 => n2220, B1 => n2221, B2 => 
                           n1880, C1 => n2222, C2 => n2192, ZN => n1720);
   U1719 : INV_X1 port map( A => n2223, ZN => n2222);
   U1720 : AND2_X1 port map( A1 => n2224, A2 => n2223, ZN => n2221);
   U1721 : OAI21_X1 port map( B1 => n2198, B2 => n2225, A => n2199, ZN => n2224
                           );
   U1722 : NAND3_X1 port map( A1 => n2195, A2 => n2223, A3 => n2226, ZN => 
                           n2220);
   U1723 : OAI21_X1 port map( B1 => n2227, B2 => n2228, A => n2181, ZN => n2223
                           );
   U1724 : OAI222_X1 port map( A1 => n2158, A2 => n2229, B1 => n2230, B2 => 
                           n1800, C1 => n2231, C2 => n2185, ZN => n1719);
   U1725 : OAI222_X1 port map( A1 => n2159, A2 => n2229, B1 => n2230, B2 => 
                           n1801, C1 => n2231, C2 => n2186, ZN => n1718);
   U1726 : OAI222_X1 port map( A1 => n2160, A2 => n2229, B1 => n2230, B2 => 
                           n1802, C1 => n2231, C2 => n2187, ZN => n1717);
   U1727 : OAI222_X1 port map( A1 => n2161, A2 => n2229, B1 => n2230, B2 => 
                           n1803, C1 => n2231, C2 => n2188, ZN => n1716);
   U1728 : OAI222_X1 port map( A1 => n2162, A2 => n2229, B1 => n2230, B2 => 
                           n1804, C1 => n2231, C2 => n2189, ZN => n1715);
   U1729 : OAI222_X1 port map( A1 => n2163, A2 => n2229, B1 => n2230, B2 => 
                           n1805, C1 => n2231, C2 => n2190, ZN => n1714);
   U1730 : OAI222_X1 port map( A1 => n2164, A2 => n2229, B1 => n2230, B2 => 
                           n1806, C1 => n2231, C2 => n2191, ZN => n1713);
   U1731 : OAI222_X1 port map( A1 => n2165, A2 => n2229, B1 => n2230, B2 => 
                           n1890, C1 => n2231, C2 => n2192, ZN => n1712);
   U1732 : INV_X1 port map( A => n2232, ZN => n2231);
   U1733 : AND2_X1 port map( A1 => n2233, A2 => n2232, ZN => n2230);
   U1734 : OAI21_X1 port map( B1 => n2198, B2 => n2234, A => n2199, ZN => n2233
                           );
   U1735 : NAND3_X1 port map( A1 => n2195, A2 => n2232, A3 => n2235, ZN => 
                           n2229);
   U1736 : OAI21_X1 port map( B1 => n2113, B2 => n2227, A => n2181, ZN => n2232
                           );
   U1737 : OAI222_X1 port map( A1 => n2158, A2 => n2236, B1 => n2237, B2 => 
                           n1953, C1 => n2238, C2 => n2185, ZN => n1711);
   U1738 : OAI222_X1 port map( A1 => n2159, A2 => n2236, B1 => n2237, B2 => 
                           n1955, C1 => n2238, C2 => n2186, ZN => n1710);
   U1739 : OAI222_X1 port map( A1 => n2160, A2 => n2236, B1 => n2237, B2 => 
                           n1957, C1 => n2238, C2 => n2187, ZN => n1709);
   U1740 : OAI222_X1 port map( A1 => n2161, A2 => n2236, B1 => n2237, B2 => 
                           n1959, C1 => n2238, C2 => n2188, ZN => n1708);
   U1741 : OAI222_X1 port map( A1 => n2162, A2 => n2236, B1 => n2237, B2 => 
                           n1961, C1 => n2238, C2 => n2189, ZN => n1707);
   U1742 : OAI222_X1 port map( A1 => n2163, A2 => n2236, B1 => n2237, B2 => 
                           n1963, C1 => n2238, C2 => n2190, ZN => n1706);
   U1743 : OAI222_X1 port map( A1 => n2164, A2 => n2236, B1 => n2237, B2 => 
                           n1965, C1 => n2238, C2 => n2191, ZN => n1705);
   U1744 : OAI222_X1 port map( A1 => n2165, A2 => n2236, B1 => n2237, B2 => 
                           n1848, C1 => n2238, C2 => n2192, ZN => n1704);
   U1745 : INV_X1 port map( A => n2239, ZN => n2238);
   U1746 : AND2_X1 port map( A1 => n2240, A2 => n2239, ZN => n2237);
   U1747 : OAI21_X1 port map( B1 => n2198, B2 => n2241, A => n2199, ZN => n2240
                           );
   U1748 : NAND3_X1 port map( A1 => n2195, A2 => n2239, A3 => n2242, ZN => 
                           n2236);
   U1749 : OAI21_X1 port map( B1 => n2227, B2 => n2243, A => n2181, ZN => n2239
                           );
   U1750 : OAI222_X1 port map( A1 => n2158, A2 => n2244, B1 => n2245, B2 => 
                           n1850, C1 => n2246, C2 => n2185, ZN => n1703);
   U1751 : OAI222_X1 port map( A1 => n2159, A2 => n2244, B1 => n2245, B2 => 
                           n1852, C1 => n2246, C2 => n2186, ZN => n1702);
   U1752 : OAI222_X1 port map( A1 => n2160, A2 => n2244, B1 => n2245, B2 => 
                           n1854, C1 => n2246, C2 => n2187, ZN => n1701);
   U1753 : OAI222_X1 port map( A1 => n2161, A2 => n2244, B1 => n2245, B2 => 
                           n1856, C1 => n2246, C2 => n2188, ZN => n1700);
   U1754 : OAI222_X1 port map( A1 => n2162, A2 => n2244, B1 => n2245, B2 => 
                           n1858, C1 => n2246, C2 => n2189, ZN => n1699);
   U1755 : OAI222_X1 port map( A1 => n2163, A2 => n2244, B1 => n2245, B2 => 
                           n1860, C1 => n2246, C2 => n2190, ZN => n1698);
   U1756 : OAI222_X1 port map( A1 => n2164, A2 => n2244, B1 => n2245, B2 => 
                           n1862, C1 => n2246, C2 => n2191, ZN => n1697);
   U1757 : OAI222_X1 port map( A1 => n2165, A2 => n2244, B1 => n2245, B2 => 
                           n1872, C1 => n2246, C2 => n2192, ZN => n1696);
   U1758 : INV_X1 port map( A => n2247, ZN => n2246);
   U1759 : AND2_X1 port map( A1 => n2248, A2 => n2247, ZN => n2245);
   U1760 : OAI21_X1 port map( B1 => n2198, B2 => n2249, A => n2199, ZN => n2248
                           );
   U1761 : NAND3_X1 port map( A1 => n2195, A2 => n2247, A3 => n2250, ZN => 
                           n2244);
   U1762 : OAI21_X1 port map( B1 => n2227, B2 => n2251, A => n2181, ZN => n2247
                           );
   U1763 : OAI222_X1 port map( A1 => n2158, A2 => n2252, B1 => n2253, B2 => 
                           n1966, C1 => n2254, C2 => n2185, ZN => n1695);
   U1764 : OAI222_X1 port map( A1 => n2159, A2 => n2252, B1 => n2253, B2 => 
                           n1967, C1 => n2254, C2 => n2186, ZN => n1694);
   U1765 : OAI222_X1 port map( A1 => n2160, A2 => n2252, B1 => n2253, B2 => 
                           n1968, C1 => n2254, C2 => n2187, ZN => n1693);
   U1766 : OAI222_X1 port map( A1 => n2161, A2 => n2252, B1 => n2253, B2 => 
                           n1969, C1 => n2254, C2 => n2188, ZN => n1692);
   U1767 : OAI222_X1 port map( A1 => n2162, A2 => n2252, B1 => n2253, B2 => 
                           n1970, C1 => n2254, C2 => n2189, ZN => n1691);
   U1768 : OAI222_X1 port map( A1 => n2163, A2 => n2252, B1 => n2253, B2 => 
                           n1971, C1 => n2254, C2 => n2190, ZN => n1690);
   U1769 : OAI222_X1 port map( A1 => n2164, A2 => n2252, B1 => n2253, B2 => 
                           n1972, C1 => n2254, C2 => n2191, ZN => n1689);
   U1770 : OAI222_X1 port map( A1 => n2165, A2 => n2252, B1 => n2253, B2 => 
                           n1996, C1 => n2254, C2 => n2192, ZN => n1688);
   U1771 : INV_X1 port map( A => n2255, ZN => n2254);
   U1772 : AND2_X1 port map( A1 => n2256, A2 => n2255, ZN => n2253);
   U1773 : OAI21_X1 port map( B1 => n2198, B2 => n2257, A => n2199, ZN => n2256
                           );
   U1774 : NAND3_X1 port map( A1 => N1665, A2 => n2180, A3 => N1666, ZN => 
                           n2198);
   U1775 : NAND3_X1 port map( A1 => n2195, A2 => n2255, A3 => n2258, ZN => 
                           n2252);
   U1776 : OAI21_X1 port map( B1 => n2115, B2 => n2227, A => n2181, ZN => n2255
                           );
   U1777 : NAND2_X1 port map( A1 => n2259, A2 => n2128, ZN => n2227);
   U1778 : AND3_X1 port map( A1 => N1666, A2 => N1665, A3 => n2260, ZN => n2195
                           );
   U1779 : OAI222_X1 port map( A1 => n2158, A2 => n2261, B1 => n2262, B2 => 
                           n1925, C1 => n2263, C2 => n2185, ZN => n1687);
   U1780 : OAI222_X1 port map( A1 => n2159, A2 => n2261, B1 => n2262, B2 => 
                           n1926, C1 => n2263, C2 => n2186, ZN => n1686);
   U1781 : OAI222_X1 port map( A1 => n2160, A2 => n2261, B1 => n2262, B2 => 
                           n1927, C1 => n2263, C2 => n2187, ZN => n1685);
   U1782 : OAI222_X1 port map( A1 => n2161, A2 => n2261, B1 => n2262, B2 => 
                           n1928, C1 => n2263, C2 => n2188, ZN => n1684);
   U1783 : OAI222_X1 port map( A1 => n2162, A2 => n2261, B1 => n2262, B2 => 
                           n1929, C1 => n2263, C2 => n2189, ZN => n1683);
   U1784 : OAI222_X1 port map( A1 => n2163, A2 => n2261, B1 => n2262, B2 => 
                           n1930, C1 => n2263, C2 => n2190, ZN => n1682);
   U1785 : OAI222_X1 port map( A1 => n2164, A2 => n2261, B1 => n2262, B2 => 
                           n1931, C1 => n2263, C2 => n2191, ZN => n1681);
   U1786 : OAI222_X1 port map( A1 => n2165, A2 => n2261, B1 => n2262, B2 => 
                           n1839, C1 => n2263, C2 => n2192, ZN => n1680);
   U1787 : INV_X1 port map( A => n2264, ZN => n2263);
   U1788 : AND2_X1 port map( A1 => n2265, A2 => n2264, ZN => n2262);
   U1789 : OAI21_X1 port map( B1 => n2197, B2 => n2266, A => n2199, ZN => n2265
                           );
   U1790 : NAND3_X1 port map( A1 => n2194, A2 => n2264, A3 => n2267, ZN => 
                           n2261);
   U1791 : OAI21_X1 port map( B1 => n2120, B2 => n2268, A => n2181, ZN => n2264
                           );
   U1792 : OAI222_X1 port map( A1 => n2158, A2 => n2269, B1 => n2270, B2 => 
                           n2006, C1 => n2271, C2 => n2185, ZN => n1679);
   U1793 : OAI222_X1 port map( A1 => n2159, A2 => n2269, B1 => n2270, B2 => 
                           n2007, C1 => n2271, C2 => n2186, ZN => n1678);
   U1794 : OAI222_X1 port map( A1 => n2160, A2 => n2269, B1 => n2270, B2 => 
                           n2008, C1 => n2271, C2 => n2187, ZN => n1677);
   U1795 : OAI222_X1 port map( A1 => n2161, A2 => n2269, B1 => n2270, B2 => 
                           n2009, C1 => n2271, C2 => n2188, ZN => n1676);
   U1796 : OAI222_X1 port map( A1 => n2162, A2 => n2269, B1 => n2270, B2 => 
                           n2010, C1 => n2271, C2 => n2189, ZN => n1675);
   U1797 : OAI222_X1 port map( A1 => n2163, A2 => n2269, B1 => n2270, B2 => 
                           n2011, C1 => n2271, C2 => n2190, ZN => n1674);
   U1798 : OAI222_X1 port map( A1 => n2164, A2 => n2269, B1 => n2270, B2 => 
                           n2012, C1 => n2271, C2 => n2191, ZN => n1673);
   U1799 : OAI222_X1 port map( A1 => n2165, A2 => n2269, B1 => n2270, B2 => 
                           n1909, C1 => n2271, C2 => n2192, ZN => n1672);
   U1800 : INV_X1 port map( A => n2272, ZN => n2271);
   U1801 : AND2_X1 port map( A1 => n2273, A2 => n2272, ZN => n2270);
   U1802 : OAI21_X1 port map( B1 => n2208, B2 => n2266, A => n2199, ZN => n2273
                           );
   U1803 : NAND3_X1 port map( A1 => n2209, A2 => n2272, A3 => n2267, ZN => 
                           n2269);
   U1804 : OAI21_X1 port map( B1 => n2274, B2 => n2268, A => n2181, ZN => n2272
                           );
   U1805 : OAI222_X1 port map( A1 => n2158, A2 => n2275, B1 => n2276, B2 => 
                           n1911, C1 => n2277, C2 => n2185, ZN => n1671);
   U1806 : OAI222_X1 port map( A1 => n2159, A2 => n2275, B1 => n2276, B2 => 
                           n1912, C1 => n2277, C2 => n2186, ZN => n1670);
   U1807 : OAI222_X1 port map( A1 => n2160, A2 => n2275, B1 => n2276, B2 => 
                           n1913, C1 => n2277, C2 => n2187, ZN => n1669);
   U1808 : OAI222_X1 port map( A1 => n2161, A2 => n2275, B1 => n2276, B2 => 
                           n1914, C1 => n2277, C2 => n2188, ZN => n1668);
   U1809 : OAI222_X1 port map( A1 => n2162, A2 => n2275, B1 => n2276, B2 => 
                           n1915, C1 => n2277, C2 => n2189, ZN => n1667);
   U1810 : OAI222_X1 port map( A1 => n2163, A2 => n2275, B1 => n2276, B2 => 
                           n1916, C1 => n2277, C2 => n2190, ZN => n1666_port);
   U1811 : OAI222_X1 port map( A1 => n2164, A2 => n2275, B1 => n2276, B2 => 
                           n1917, C1 => n2277, C2 => n2191, ZN => n1665_port);
   U1812 : OAI222_X1 port map( A1 => n2165, A2 => n2275, B1 => n2276, B2 => 
                           n1871, C1 => n2277, C2 => n2192, ZN => n1664_port);
   U1813 : INV_X1 port map( A => n2278, ZN => n2277);
   U1814 : AND2_X1 port map( A1 => n2279, A2 => n2278, ZN => n2276);
   U1815 : OAI21_X1 port map( B1 => n2216, B2 => n2266, A => n2199, ZN => n2279
                           );
   U1816 : NAND3_X1 port map( A1 => n2217, A2 => n2278, A3 => n2267, ZN => 
                           n2275);
   U1817 : OAI21_X1 port map( B1 => n2219, B2 => n2280, A => n2181, ZN => n2278
                           );
   U1818 : OAI222_X1 port map( A1 => n2158, A2 => n2281, B1 => n2282, B2 => 
                           n1988, C1 => n2283, C2 => n2185, ZN => n1663_port);
   U1819 : INV_X1 port map( A => DATAIN(0), ZN => n2158);
   U1820 : OAI222_X1 port map( A1 => n2159, A2 => n2281, B1 => n2282, B2 => 
                           n1989, C1 => n2283, C2 => n2186, ZN => n1662_port);
   U1821 : INV_X1 port map( A => DATAIN(1), ZN => n2159);
   U1822 : OAI222_X1 port map( A1 => n2160, A2 => n2281, B1 => n2282, B2 => 
                           n1990, C1 => n2283, C2 => n2187, ZN => n1661);
   U1823 : INV_X1 port map( A => DATAIN(2), ZN => n2160);
   U1824 : OAI222_X1 port map( A1 => n2161, A2 => n2281, B1 => n2282, B2 => 
                           n1991, C1 => n2283, C2 => n2188, ZN => n1660);
   U1825 : INV_X1 port map( A => DATAIN(3), ZN => n2161);
   U1826 : OAI222_X1 port map( A1 => n2162, A2 => n2281, B1 => n2282, B2 => 
                           n1992, C1 => n2283, C2 => n2189, ZN => n1659);
   U1827 : INV_X1 port map( A => DATAIN(4), ZN => n2162);
   U1828 : OAI222_X1 port map( A1 => n2163, A2 => n2281, B1 => n2282, B2 => 
                           n1993, C1 => n2283, C2 => n2190, ZN => n1658);
   U1829 : INV_X1 port map( A => DATAIN(5), ZN => n2163);
   U1830 : OAI222_X1 port map( A1 => n2164, A2 => n2281, B1 => n2282, B2 => 
                           n1994, C1 => n2283, C2 => n2191, ZN => n1657);
   U1831 : INV_X1 port map( A => DATAIN(6), ZN => n2164);
   U1832 : OAI222_X1 port map( A1 => n2165, A2 => n2281, B1 => n2282, B2 => 
                           n1995, C1 => n2283, C2 => n2192, ZN => n1656);
   U1833 : INV_X1 port map( A => n2284, ZN => n2283);
   U1834 : AND2_X1 port map( A1 => n2285, A2 => n2284, ZN => n2282);
   U1835 : OAI21_X1 port map( B1 => n2225, B2 => n2266, A => n2199, ZN => n2285
                           );
   U1836 : NAND2_X1 port map( A1 => n2286, A2 => n2180, ZN => n2266);
   U1837 : NAND3_X1 port map( A1 => n2226, A2 => n2284, A3 => n2267, ZN => 
                           n2281);
   U1838 : AND2_X1 port map( A1 => n2286, A2 => n2260, ZN => n2267);
   U1839 : OAI21_X1 port map( B1 => n2219, B2 => n2287, A => n2181, ZN => n2284
                           );
   U1840 : INV_X1 port map( A => DATAIN(7), ZN => n2165);
   U1841 : OAI222_X1 port map( A1 => n2288, A2 => n1873, B1 => n2289, B2 => 
                           n2290, C1 => n2185, C2 => n2291, ZN => n1655);
   U1842 : OAI222_X1 port map( A1 => n2288, A2 => n1874, B1 => n2289, B2 => 
                           n2292, C1 => n2186, C2 => n2291, ZN => n1654);
   U1843 : OAI222_X1 port map( A1 => n2288, A2 => n1875, B1 => n2289, B2 => 
                           n2293, C1 => n2187, C2 => n2291, ZN => n1653);
   U1844 : OAI222_X1 port map( A1 => n2288, A2 => n1876, B1 => n2289, B2 => 
                           n2294, C1 => n2188, C2 => n2291, ZN => n1652);
   U1845 : OAI222_X1 port map( A1 => n2288, A2 => n1877, B1 => n2289, B2 => 
                           n2295, C1 => n2189, C2 => n2291, ZN => n1651);
   U1846 : OAI222_X1 port map( A1 => n2288, A2 => n1878, B1 => n2289, B2 => 
                           n2296, C1 => n2190, C2 => n2291, ZN => n1650);
   U1847 : OAI222_X1 port map( A1 => n2288, A2 => n1879, B1 => n2289, B2 => 
                           n2297, C1 => n2191, C2 => n2291, ZN => n1649);
   U1848 : OAI222_X1 port map( A1 => n2288, A2 => n1815, B1 => n2289, B2 => 
                           n2298, C1 => n2192, C2 => n2291, ZN => n1648);
   U1849 : NAND3_X1 port map( A1 => n2286, A2 => n2235, A3 => n2299, ZN => 
                           n2289);
   U1850 : AND3_X1 port map( A1 => n2299, A2 => n2300, A3 => n2301, ZN => n2288
                           );
   U1851 : INV_X1 port map( A => n2291, ZN => n2299);
   U1852 : OAI21_X1 port map( B1 => n2302, B2 => n2201, A => n2202, ZN => n2291
                           );
   U1853 : OAI222_X1 port map( A1 => n2290, A2 => n2303, B1 => n2304, B2 => 
                           n2013, C1 => n2305, C2 => n2185, ZN => n1647);
   U1854 : OAI222_X1 port map( A1 => n2292, A2 => n2303, B1 => n2304, B2 => 
                           n2014, C1 => n2305, C2 => n2186, ZN => n1646);
   U1855 : OAI222_X1 port map( A1 => n2293, A2 => n2303, B1 => n2304, B2 => 
                           n2015, C1 => n2305, C2 => n2187, ZN => n1645);
   U1856 : OAI222_X1 port map( A1 => n2294, A2 => n2303, B1 => n2304, B2 => 
                           n2016, C1 => n2305, C2 => n2188, ZN => n1644);
   U1857 : OAI222_X1 port map( A1 => n2295, A2 => n2303, B1 => n2304, B2 => 
                           n2017, C1 => n2305, C2 => n2189, ZN => n1643);
   U1858 : OAI222_X1 port map( A1 => n2296, A2 => n2303, B1 => n2304, B2 => 
                           n2018, C1 => n2305, C2 => n2190, ZN => n1642);
   U1859 : OAI222_X1 port map( A1 => n2297, A2 => n2303, B1 => n2304, B2 => 
                           n2019, C1 => n2305, C2 => n2191, ZN => n1641);
   U1860 : OAI222_X1 port map( A1 => n2298, A2 => n2303, B1 => n2304, B2 => 
                           n1908, C1 => n2305, C2 => n2192, ZN => n1640);
   U1861 : INV_X1 port map( A => n2306, ZN => n2305);
   U1862 : AND3_X1 port map( A1 => n2307, A2 => n2306, A3 => n2301, ZN => n2304
                           );
   U1863 : NAND3_X1 port map( A1 => n2242, A2 => n2306, A3 => n2286, ZN => 
                           n2303);
   U1864 : OAI21_X1 port map( B1 => n2243, B2 => n2268, A => n2181, ZN => n2306
                           );
   U1865 : OAI222_X1 port map( A1 => n2290, A2 => n2308, B1 => n2309, B2 => 
                           n1973, C1 => n2185, C2 => n2310, ZN => n1639);
   U1866 : OAI222_X1 port map( A1 => n2292, A2 => n2308, B1 => n2309, B2 => 
                           n1974, C1 => n2186, C2 => n2310, ZN => n1638);
   U1867 : OAI222_X1 port map( A1 => n2293, A2 => n2308, B1 => n2309, B2 => 
                           n1975, C1 => n2187, C2 => n2310, ZN => n1637);
   U1868 : OAI222_X1 port map( A1 => n2294, A2 => n2308, B1 => n2309, B2 => 
                           n1976, C1 => n2188, C2 => n2310, ZN => n1636);
   U1869 : OAI222_X1 port map( A1 => n2295, A2 => n2308, B1 => n2309, B2 => 
                           n1977, C1 => n2189, C2 => n2310, ZN => n1635);
   U1870 : OAI222_X1 port map( A1 => n2296, A2 => n2308, B1 => n2309, B2 => 
                           n1978, C1 => n2190, C2 => n2310, ZN => n1634);
   U1871 : OAI222_X1 port map( A1 => n2297, A2 => n2308, B1 => n2309, B2 => 
                           n1979, C1 => n2191, C2 => n2310, ZN => n1633);
   U1872 : OAI222_X1 port map( A1 => n2298, A2 => n2308, B1 => n2309, B2 => 
                           n1980, C1 => n2192, C2 => n2310, ZN => n1632);
   U1873 : AND3_X1 port map( A1 => n2301, A2 => n2311, A3 => n2312, ZN => n2309
                           );
   U1874 : NAND3_X1 port map( A1 => n2286, A2 => n2250, A3 => n2312, ZN => 
                           n2308);
   U1875 : INV_X1 port map( A => n2310, ZN => n2312);
   U1876 : OAI21_X1 port map( B1 => n2313, B2 => n2201, A => n2202, ZN => n2310
                           );
   U1877 : OAI222_X1 port map( A1 => n2290, A2 => n2314, B1 => n2315, B2 => 
                           n2020, C1 => n2316, C2 => n2185, ZN => n1631);
   U1878 : OAI222_X1 port map( A1 => n2292, A2 => n2314, B1 => n2315, B2 => 
                           n2021, C1 => n2316, C2 => n2186, ZN => n1630);
   U1879 : OAI222_X1 port map( A1 => n2293, A2 => n2314, B1 => n2315, B2 => 
                           n2022, C1 => n2316, C2 => n2187, ZN => n1629);
   U1880 : OAI222_X1 port map( A1 => n2294, A2 => n2314, B1 => n2315, B2 => 
                           n2023, C1 => n2316, C2 => n2188, ZN => n1628);
   U1881 : OAI222_X1 port map( A1 => n2295, A2 => n2314, B1 => n2315, B2 => 
                           n2024, C1 => n2316, C2 => n2189, ZN => n1627);
   U1882 : OAI222_X1 port map( A1 => n2296, A2 => n2314, B1 => n2315, B2 => 
                           n2025, C1 => n2316, C2 => n2190, ZN => n1626);
   U1883 : OAI222_X1 port map( A1 => n2297, A2 => n2314, B1 => n2315, B2 => 
                           n2026, C1 => n2316, C2 => n2191, ZN => n1625);
   U1884 : OAI222_X1 port map( A1 => n2298, A2 => n2314, B1 => n2315, B2 => 
                           n2027, C1 => n2316, C2 => n2192, ZN => n1624);
   U1885 : INV_X1 port map( A => n2317, ZN => n2316);
   U1886 : AND3_X1 port map( A1 => n2318, A2 => n2317, A3 => n2301, ZN => n2315
                           );
   U1887 : INV_X1 port map( A => n2319, ZN => n2301);
   U1888 : OAI21_X1 port map( B1 => n2286, B2 => n2132, A => n2320, ZN => n2319
                           );
   U1889 : NAND3_X1 port map( A1 => n2258, A2 => n2317, A3 => n2286, ZN => 
                           n2314);
   U1890 : NOR2_X1 port map( A1 => n2151, A2 => N1665, ZN => n2286);
   U1891 : INV_X1 port map( A => N1666, ZN => n2151);
   U1892 : OAI21_X1 port map( B1 => n2115, B2 => n2268, A => n2181, ZN => n2317
                           );
   U1893 : NAND2_X1 port map( A1 => n2125, A2 => n2259, ZN => n2268);
   U1894 : OAI222_X1 port map( A1 => n2290, A2 => n2321, B1 => n3191, B2 => 
                           n2322, C1 => n2323, C2 => n2185, ZN => n1623);
   U1895 : OAI222_X1 port map( A1 => n2292, A2 => n2321, B1 => n3179, B2 => 
                           n2322, C1 => n2323, C2 => n2186, ZN => n1622);
   U1896 : OAI222_X1 port map( A1 => n2293, A2 => n2321, B1 => n3167, B2 => 
                           n2322, C1 => n2323, C2 => n2187, ZN => n1621);
   U1897 : OAI222_X1 port map( A1 => n2294, A2 => n2321, B1 => n3155, B2 => 
                           n2322, C1 => n2323, C2 => n2188, ZN => n1620);
   U1898 : OAI222_X1 port map( A1 => n2295, A2 => n2321, B1 => n3143, B2 => 
                           n2322, C1 => n2323, C2 => n2189, ZN => n1619);
   U1899 : OAI222_X1 port map( A1 => n2296, A2 => n2321, B1 => n3131, B2 => 
                           n2322, C1 => n2323, C2 => n2190, ZN => n1618);
   U1900 : OAI222_X1 port map( A1 => n2297, A2 => n2321, B1 => n3119, B2 => 
                           n2322, C1 => n2323, C2 => n2191, ZN => n1617);
   U1901 : OAI222_X1 port map( A1 => n2298, A2 => n2321, B1 => n3109, B2 => 
                           n2322, C1 => n2323, C2 => n2192, ZN => n1616);
   U1902 : INV_X1 port map( A => n2324, ZN => n2323);
   U1903 : AND3_X1 port map( A1 => n2325, A2 => n2324, A3 => n2326, ZN => n2322
                           );
   U1904 : NAND3_X1 port map( A1 => n2194, A2 => n2324, A3 => n2327, ZN => 
                           n2321);
   U1905 : OAI21_X1 port map( B1 => n2219, B2 => n2126, A => n2181, ZN => n2324
                           );
   U1906 : OAI222_X1 port map( A1 => n2290, A2 => n2328, B1 => n2329, B2 => 
                           n1981, C1 => n2330, C2 => n2185, ZN => n1615);
   U1907 : OAI222_X1 port map( A1 => n2292, A2 => n2328, B1 => n2329, B2 => 
                           n1982, C1 => n2330, C2 => n2186, ZN => n1614);
   U1908 : OAI222_X1 port map( A1 => n2293, A2 => n2328, B1 => n2329, B2 => 
                           n1983, C1 => n2330, C2 => n2187, ZN => n1613);
   U1909 : OAI222_X1 port map( A1 => n2294, A2 => n2328, B1 => n2329, B2 => 
                           n1984, C1 => n2330, C2 => n2188, ZN => n1612);
   U1910 : OAI222_X1 port map( A1 => n2295, A2 => n2328, B1 => n2329, B2 => 
                           n1985, C1 => n2330, C2 => n2189, ZN => n1611);
   U1911 : OAI222_X1 port map( A1 => n2296, A2 => n2328, B1 => n2329, B2 => 
                           n1986, C1 => n2330, C2 => n2190, ZN => n1610);
   U1912 : OAI222_X1 port map( A1 => n2297, A2 => n2328, B1 => n2329, B2 => 
                           n1987, C1 => n2330, C2 => n2191, ZN => n1609);
   U1913 : OAI222_X1 port map( A1 => n2298, A2 => n2328, B1 => n2329, B2 => 
                           n1799, C1 => n2330, C2 => n2192, ZN => n1608);
   U1914 : INV_X1 port map( A => n2331, ZN => n2330);
   U1915 : AND3_X1 port map( A1 => n2332, A2 => n2331, A3 => n2326, ZN => n2329
                           );
   U1916 : NAND3_X1 port map( A1 => n2209, A2 => n2331, A3 => n2327, ZN => 
                           n2328);
   U1917 : OAI21_X1 port map( B1 => n2274, B2 => n2333, A => n2181, ZN => n2331
                           );
   U1918 : OAI222_X1 port map( A1 => n2290, A2 => n2334, B1 => n3029, B2 => 
                           n2335, C1 => n2336, C2 => n2185, ZN => n1607);
   U1919 : OAI222_X1 port map( A1 => n2292, A2 => n2334, B1 => n3030, B2 => 
                           n2335, C1 => n2336, C2 => n2186, ZN => n1606);
   U1920 : OAI222_X1 port map( A1 => n2293, A2 => n2334, B1 => n3031, B2 => 
                           n2335, C1 => n2336, C2 => n2187, ZN => n1605);
   U1921 : OAI222_X1 port map( A1 => n2294, A2 => n2334, B1 => n3032, B2 => 
                           n2335, C1 => n2336, C2 => n2188, ZN => n1604);
   U1922 : OAI222_X1 port map( A1 => n2295, A2 => n2334, B1 => n3033, B2 => 
                           n2335, C1 => n2336, C2 => n2189, ZN => n1603);
   U1923 : OAI222_X1 port map( A1 => n2296, A2 => n2334, B1 => n3034, B2 => 
                           n2335, C1 => n2336, C2 => n2190, ZN => n1602);
   U1924 : OAI222_X1 port map( A1 => n2297, A2 => n2334, B1 => n3035, B2 => 
                           n2335, C1 => n2336, C2 => n2191, ZN => n1601);
   U1925 : OAI222_X1 port map( A1 => n2298, A2 => n2334, B1 => n3036, B2 => 
                           n2335, C1 => n2336, C2 => n2192, ZN => n1600);
   U1926 : INV_X1 port map( A => n2337, ZN => n2336);
   U1927 : AND3_X1 port map( A1 => n2338, A2 => n2337, A3 => n2326, ZN => n2335
                           );
   U1928 : NAND3_X1 port map( A1 => n2217, A2 => n2337, A3 => n2327, ZN => 
                           n2334);
   U1929 : OAI21_X1 port map( B1 => n2339, B2 => n2333, A => n2181, ZN => n2337
                           );
   U1930 : OAI222_X1 port map( A1 => n2290, A2 => n2340, B1 => n3274, B2 => 
                           n2341, C1 => n2342, C2 => n2185, ZN => n1599);
   U1931 : OAI222_X1 port map( A1 => n2292, A2 => n2340, B1 => n3266, B2 => 
                           n2341, C1 => n2342, C2 => n2186, ZN => n1598);
   U1932 : OAI222_X1 port map( A1 => n2293, A2 => n2340, B1 => n3258, B2 => 
                           n2341, C1 => n2342, C2 => n2187, ZN => n1597);
   U1933 : OAI222_X1 port map( A1 => n2294, A2 => n2340, B1 => n3250, B2 => 
                           n2341, C1 => n2342, C2 => n2188, ZN => n1596);
   U1934 : OAI222_X1 port map( A1 => n2295, A2 => n2340, B1 => n3242, B2 => 
                           n2341, C1 => n2342, C2 => n2189, ZN => n1595);
   U1935 : OAI222_X1 port map( A1 => n2296, A2 => n2340, B1 => n3234, B2 => 
                           n2341, C1 => n2342, C2 => n2190, ZN => n1594);
   U1936 : OAI222_X1 port map( A1 => n2297, A2 => n2340, B1 => n3226, B2 => 
                           n2341, C1 => n2342, C2 => n2191, ZN => n1593);
   U1937 : OAI222_X1 port map( A1 => n2298, A2 => n2340, B1 => n3220, B2 => 
                           n2341, C1 => n2342, C2 => n2192, ZN => n1592);
   U1938 : INV_X1 port map( A => n2343, ZN => n2342);
   U1939 : AND3_X1 port map( A1 => n2344, A2 => n2343, A3 => n2326, ZN => n2341
                           );
   U1940 : NAND3_X1 port map( A1 => n2226, A2 => n2343, A3 => n2327, ZN => 
                           n2340);
   U1941 : OAI21_X1 port map( B1 => n2219, B2 => n2345, A => n2181, ZN => n2343
                           );
   U1942 : OAI222_X1 port map( A1 => n2290, A2 => n2346, B1 => n2347, B2 => 
                           n1831, C1 => n2348, C2 => n2185, ZN => n1591);
   U1943 : OAI222_X1 port map( A1 => n2292, A2 => n2346, B1 => n2347, B2 => 
                           n1832, C1 => n2348, C2 => n2186, ZN => n1590);
   U1944 : OAI222_X1 port map( A1 => n2293, A2 => n2346, B1 => n2347, B2 => 
                           n1833, C1 => n2348, C2 => n2187, ZN => n1589);
   U1945 : OAI222_X1 port map( A1 => n2294, A2 => n2346, B1 => n2347, B2 => 
                           n1834, C1 => n2348, C2 => n2188, ZN => n1588);
   U1946 : OAI222_X1 port map( A1 => n2295, A2 => n2346, B1 => n2347, B2 => 
                           n1835, C1 => n2348, C2 => n2189, ZN => n1587);
   U1947 : OAI222_X1 port map( A1 => n2296, A2 => n2346, B1 => n2347, B2 => 
                           n1836, C1 => n2348, C2 => n2190, ZN => n1586);
   U1948 : OAI222_X1 port map( A1 => n2297, A2 => n2346, B1 => n2347, B2 => 
                           n1837, C1 => n2348, C2 => n2191, ZN => n1585);
   U1949 : OAI222_X1 port map( A1 => n2298, A2 => n2346, B1 => n2347, B2 => 
                           n1838, C1 => n2348, C2 => n2192, ZN => n1584);
   U1950 : INV_X1 port map( A => n2349, ZN => n2348);
   U1951 : AND3_X1 port map( A1 => n2349, A2 => n2300, A3 => n2326, ZN => n2347
                           );
   U1952 : NAND3_X1 port map( A1 => n2235, A2 => n2349, A3 => n2327, ZN => 
                           n2346);
   U1953 : OAI21_X1 port map( B1 => n2113, B2 => n2333, A => n2181, ZN => n2349
                           );
   U1954 : OAI222_X1 port map( A1 => n2290, A2 => n2350, B1 => n3276, B2 => 
                           n2351, C1 => n2352, C2 => n2185, ZN => n1583);
   U1955 : OAI222_X1 port map( A1 => n2292, A2 => n2350, B1 => n3268, B2 => 
                           n2351, C1 => n2352, C2 => n2186, ZN => n1582);
   U1956 : OAI222_X1 port map( A1 => n2293, A2 => n2350, B1 => n3260, B2 => 
                           n2351, C1 => n2352, C2 => n2187, ZN => n1581);
   U1957 : OAI222_X1 port map( A1 => n2294, A2 => n2350, B1 => n3252, B2 => 
                           n2351, C1 => n2352, C2 => n2188, ZN => n1580);
   U1958 : OAI222_X1 port map( A1 => n2295, A2 => n2350, B1 => n3244, B2 => 
                           n2351, C1 => n2352, C2 => n2189, ZN => n1579);
   U1959 : OAI222_X1 port map( A1 => n2296, A2 => n2350, B1 => n3236, B2 => 
                           n2351, C1 => n2352, C2 => n2190, ZN => n1578);
   U1960 : OAI222_X1 port map( A1 => n2297, A2 => n2350, B1 => n3228, B2 => 
                           n2351, C1 => n2352, C2 => n2191, ZN => n1577);
   U1961 : OAI222_X1 port map( A1 => n2298, A2 => n2350, B1 => n3222, B2 => 
                           n2351, C1 => n2352, C2 => n2192, ZN => n1576);
   U1962 : INV_X1 port map( A => n2353, ZN => n2352);
   U1963 : AND3_X1 port map( A1 => n2353, A2 => n2307, A3 => n2326, ZN => n2351
                           );
   U1964 : NAND3_X1 port map( A1 => n2242, A2 => n2353, A3 => n2327, ZN => 
                           n2350);
   U1965 : OAI21_X1 port map( B1 => n2219, B2 => n2354, A => n2181, ZN => n2353
                           );
   U1966 : OAI222_X1 port map( A1 => n2290, A2 => n2355, B1 => n2356, B2 => 
                           n1808, C1 => n2357, C2 => n2185, ZN => n1575);
   U1967 : OAI222_X1 port map( A1 => n2292, A2 => n2355, B1 => n2356, B2 => 
                           n1809, C1 => n2357, C2 => n2186, ZN => n1574);
   U1968 : OAI222_X1 port map( A1 => n2293, A2 => n2355, B1 => n2356, B2 => 
                           n1810, C1 => n2357, C2 => n2187, ZN => n1573);
   U1969 : OAI222_X1 port map( A1 => n2294, A2 => n2355, B1 => n2356, B2 => 
                           n1811, C1 => n2357, C2 => n2188, ZN => n1572);
   U1970 : OAI222_X1 port map( A1 => n2295, A2 => n2355, B1 => n2356, B2 => 
                           n1812, C1 => n2357, C2 => n2189, ZN => n1571);
   U1971 : OAI222_X1 port map( A1 => n2296, A2 => n2355, B1 => n2356, B2 => 
                           n1813, C1 => n2357, C2 => n2190, ZN => n1570);
   U1972 : OAI222_X1 port map( A1 => n2297, A2 => n2355, B1 => n2356, B2 => 
                           n1814, C1 => n2357, C2 => n2191, ZN => n1569);
   U1973 : OAI222_X1 port map( A1 => n2298, A2 => n2355, B1 => n2356, B2 => 
                           n1891, C1 => n2357, C2 => n2192, ZN => n1568);
   U1974 : INV_X1 port map( A => n2358, ZN => n2357);
   U1975 : AND3_X1 port map( A1 => n2358, A2 => n2311, A3 => n2326, ZN => n2356
                           );
   U1976 : NAND3_X1 port map( A1 => n2250, A2 => n2358, A3 => n2327, ZN => 
                           n2355);
   U1977 : OAI21_X1 port map( B1 => n2251, B2 => n2333, A => n2181, ZN => n2358
                           );
   U1978 : NAND2_X1 port map( A1 => n2259, A2 => n2359, ZN => n2333);
   U1979 : OAI222_X1 port map( A1 => n2290, A2 => n2360, B1 => n3275, B2 => 
                           n2361, C1 => n2185, C2 => n2362, ZN => n1567);
   U1980 : OAI222_X1 port map( A1 => n2292, A2 => n2360, B1 => n3267, B2 => 
                           n2361, C1 => n2186, C2 => n2362, ZN => n1566);
   U1981 : OAI222_X1 port map( A1 => n2293, A2 => n2360, B1 => n3259, B2 => 
                           n2361, C1 => n2187, C2 => n2362, ZN => n1565);
   U1982 : OAI222_X1 port map( A1 => n2294, A2 => n2360, B1 => n3251, B2 => 
                           n2361, C1 => n2188, C2 => n2362, ZN => n1564);
   U1983 : OAI222_X1 port map( A1 => n2295, A2 => n2360, B1 => n3243, B2 => 
                           n2361, C1 => n2189, C2 => n2362, ZN => n1563);
   U1984 : OAI222_X1 port map( A1 => n2296, A2 => n2360, B1 => n3235, B2 => 
                           n2361, C1 => n2190, C2 => n2362, ZN => n1562);
   U1985 : OAI222_X1 port map( A1 => n2297, A2 => n2360, B1 => n3227, B2 => 
                           n2361, C1 => n2191, C2 => n2362, ZN => n1561);
   U1986 : OAI222_X1 port map( A1 => n2298, A2 => n2360, B1 => n3221, B2 => 
                           n2361, C1 => n2192, C2 => n2362, ZN => n1560);
   U1987 : AND3_X1 port map( A1 => n2326, A2 => n2318, A3 => n2363, ZN => n2361
                           );
   U1988 : INV_X1 port map( A => n2364, ZN => n2326);
   U1989 : OAI21_X1 port map( B1 => n2327, B2 => n2132, A => n2320, ZN => n2364
                           );
   U1990 : NAND3_X1 port map( A1 => n2327, A2 => n2258, A3 => n2363, ZN => 
                           n2360);
   U1991 : INV_X1 port map( A => n2362, ZN => n2363);
   U1992 : OAI21_X1 port map( B1 => n2365, B2 => n2201, A => n2202, ZN => n2362
                           );
   U1993 : NOR2_X1 port map( A1 => n2150, A2 => N1666, ZN => n2327);
   U1994 : INV_X1 port map( A => N1665, ZN => n2150);
   U1995 : OAI222_X1 port map( A1 => n2290, A2 => n2366, B1 => n2367, B2 => 
                           n1894, C1 => n2185, C2 => n2368, ZN => n1559);
   U1996 : OAI222_X1 port map( A1 => n2292, A2 => n2366, B1 => n2367, B2 => 
                           n1895, C1 => n2186, C2 => n2368, ZN => n1558);
   U1997 : OAI222_X1 port map( A1 => n2293, A2 => n2366, B1 => n2367, B2 => 
                           n1896, C1 => n2187, C2 => n2368, ZN => n1557);
   U1998 : OAI222_X1 port map( A1 => n2294, A2 => n2366, B1 => n2367, B2 => 
                           n1897, C1 => n2188, C2 => n2368, ZN => n1556);
   U1999 : OAI222_X1 port map( A1 => n2295, A2 => n2366, B1 => n2367, B2 => 
                           n1898, C1 => n2189, C2 => n2368, ZN => n1555);
   U2000 : OAI222_X1 port map( A1 => n2296, A2 => n2366, B1 => n2367, B2 => 
                           n1899, C1 => n2190, C2 => n2368, ZN => n1554);
   U2001 : OAI222_X1 port map( A1 => n2297, A2 => n2366, B1 => n2367, B2 => 
                           n1900, C1 => n2191, C2 => n2368, ZN => n1553);
   U2002 : OAI222_X1 port map( A1 => n2298, A2 => n2366, B1 => n2367, B2 => 
                           n1901, C1 => n2192, C2 => n2368, ZN => n1552);
   U2003 : AND3_X1 port map( A1 => n2369, A2 => n2325, A3 => n2370, ZN => n2367
                           );
   U2004 : NAND2_X1 port map( A1 => n2199, A2 => n2197, ZN => n2325);
   U2005 : NAND3_X1 port map( A1 => n2370, A2 => n2194, A3 => n2371, ZN => 
                           n2366);
   U2006 : INV_X1 port map( A => n2197, ZN => n2194);
   U2007 : NAND3_X1 port map( A1 => N1663, A2 => N1662, A3 => N1664, ZN => 
                           n2197);
   U2008 : INV_X1 port map( A => n2368, ZN => n2370);
   U2009 : OAI21_X1 port map( B1 => n2372, B2 => n2201, A => n2202, ZN => n2368
                           );
   U2010 : OAI222_X1 port map( A1 => n2290, A2 => n2373, B1 => n2374, B2 => 
                           n2028, C1 => n2375, C2 => n2185, ZN => n1551);
   U2011 : OAI222_X1 port map( A1 => n2292, A2 => n2373, B1 => n2374, B2 => 
                           n2029, C1 => n2375, C2 => n2186, ZN => n1550);
   U2012 : OAI222_X1 port map( A1 => n2293, A2 => n2373, B1 => n2374, B2 => 
                           n2030, C1 => n2375, C2 => n2187, ZN => n1549);
   U2013 : OAI222_X1 port map( A1 => n2294, A2 => n2373, B1 => n2374, B2 => 
                           n2031, C1 => n2375, C2 => n2188, ZN => n1548);
   U2014 : OAI222_X1 port map( A1 => n2295, A2 => n2373, B1 => n2374, B2 => 
                           n2032, C1 => n2375, C2 => n2189, ZN => n1547);
   U2015 : OAI222_X1 port map( A1 => n2296, A2 => n2373, B1 => n2374, B2 => 
                           n2033, C1 => n2375, C2 => n2190, ZN => n1546);
   U2016 : OAI222_X1 port map( A1 => n2297, A2 => n2373, B1 => n2374, B2 => 
                           n2034, C1 => n2375, C2 => n2191, ZN => n1545);
   U2017 : OAI222_X1 port map( A1 => n2298, A2 => n2373, B1 => n2374, B2 => 
                           n1907, C1 => n2375, C2 => n2192, ZN => n1544);
   U2018 : INV_X1 port map( A => n2376, ZN => n2375);
   U2019 : AND3_X1 port map( A1 => n2376, A2 => n2332, A3 => n2369, ZN => n2374
                           );
   U2020 : NAND2_X1 port map( A1 => n2199, A2 => n2208, ZN => n2332);
   U2021 : NAND3_X1 port map( A1 => n2209, A2 => n2376, A3 => n2371, ZN => 
                           n2373);
   U2022 : OAI21_X1 port map( B1 => n2274, B2 => n2377, A => n2181, ZN => n2376
                           );
   U2023 : INV_X1 port map( A => n2208, ZN => n2209);
   U2024 : NAND3_X1 port map( A1 => N1663, A2 => n2147, A3 => N1664, ZN => 
                           n2208);
   U2025 : OAI222_X1 port map( A1 => n2290, A2 => n2378, B1 => n3196, B2 => 
                           n2379, C1 => n2380, C2 => n2185, ZN => n1543);
   U2026 : OAI222_X1 port map( A1 => n2292, A2 => n2378, B1 => n3184, B2 => 
                           n2379, C1 => n2380, C2 => n2186, ZN => n1542);
   U2027 : OAI222_X1 port map( A1 => n2293, A2 => n2378, B1 => n3172, B2 => 
                           n2379, C1 => n2380, C2 => n2187, ZN => n1541);
   U2028 : OAI222_X1 port map( A1 => n2294, A2 => n2378, B1 => n3160, B2 => 
                           n2379, C1 => n2380, C2 => n2188, ZN => n1540);
   U2029 : OAI222_X1 port map( A1 => n2295, A2 => n2378, B1 => n3148, B2 => 
                           n2379, C1 => n2380, C2 => n2189, ZN => n1539);
   U2030 : OAI222_X1 port map( A1 => n2296, A2 => n2378, B1 => n3136, B2 => 
                           n2379, C1 => n2380, C2 => n2190, ZN => n1538);
   U2031 : OAI222_X1 port map( A1 => n2297, A2 => n2378, B1 => n3124, B2 => 
                           n2379, C1 => n2380, C2 => n2191, ZN => n1537);
   U2032 : OAI222_X1 port map( A1 => n2298, A2 => n2378, B1 => n3114, B2 => 
                           n2379, C1 => n2380, C2 => n2192, ZN => n1536);
   U2033 : INV_X1 port map( A => n2381, ZN => n2380);
   U2034 : AND3_X1 port map( A1 => n2381, A2 => n2338, A3 => n2369, ZN => n2379
                           );
   U2035 : NAND2_X1 port map( A1 => n2199, A2 => n2216, ZN => n2338);
   U2036 : NAND3_X1 port map( A1 => n2217, A2 => n2381, A3 => n2371, ZN => 
                           n2378);
   U2037 : OAI21_X1 port map( B1 => n2219, B2 => n2382, A => n2181, ZN => n2381
                           );
   U2038 : INV_X1 port map( A => n2216, ZN => n2217);
   U2039 : NAND3_X1 port map( A1 => N1662, A2 => n2148, A3 => N1664, ZN => 
                           n2216);
   U2040 : OAI222_X1 port map( A1 => n2290, A2 => n2383, B1 => n2384, B2 => 
                           n1823, C1 => n2385, C2 => n2185, ZN => n1535);
   U2041 : OAI222_X1 port map( A1 => n2292, A2 => n2383, B1 => n2384, B2 => 
                           n1824, C1 => n2385, C2 => n2186, ZN => n1534);
   U2042 : OAI222_X1 port map( A1 => n2293, A2 => n2383, B1 => n2384, B2 => 
                           n1825, C1 => n2385, C2 => n2187, ZN => n1533);
   U2043 : OAI222_X1 port map( A1 => n2294, A2 => n2383, B1 => n2384, B2 => 
                           n1826, C1 => n2385, C2 => n2188, ZN => n1532);
   U2044 : OAI222_X1 port map( A1 => n2295, A2 => n2383, B1 => n2384, B2 => 
                           n1827, C1 => n2385, C2 => n2189, ZN => n1531);
   U2045 : OAI222_X1 port map( A1 => n2296, A2 => n2383, B1 => n2384, B2 => 
                           n1828, C1 => n2385, C2 => n2190, ZN => n1530);
   U2046 : OAI222_X1 port map( A1 => n2297, A2 => n2383, B1 => n2384, B2 => 
                           n1829, C1 => n2385, C2 => n2191, ZN => n1529);
   U2047 : OAI222_X1 port map( A1 => n2298, A2 => n2383, B1 => n2384, B2 => 
                           n1881, C1 => n2385, C2 => n2192, ZN => n1528);
   U2048 : INV_X1 port map( A => n2386, ZN => n2385);
   U2049 : AND3_X1 port map( A1 => n2386, A2 => n2344, A3 => n2369, ZN => n2384
                           );
   U2050 : NAND2_X1 port map( A1 => n2199, A2 => n2225, ZN => n2344);
   U2051 : NAND3_X1 port map( A1 => n2226, A2 => n2386, A3 => n2371, ZN => 
                           n2383);
   U2052 : OAI21_X1 port map( B1 => n2228, B2 => n2377, A => n2181, ZN => n2386
                           );
   U2053 : INV_X1 port map( A => n2225, ZN => n2226);
   U2054 : NAND3_X1 port map( A1 => n2147, A2 => n2148, A3 => N1664, ZN => 
                           n2225);
   U2055 : OAI222_X1 port map( A1 => n2290, A2 => n2387, B1 => n3194, B2 => 
                           n2388, C1 => n2389, C2 => n2185, ZN => n1527);
   U2056 : OAI222_X1 port map( A1 => n2292, A2 => n2387, B1 => n3182, B2 => 
                           n2388, C1 => n2389, C2 => n2186, ZN => n1526);
   U2057 : OAI222_X1 port map( A1 => n2293, A2 => n2387, B1 => n3170, B2 => 
                           n2388, C1 => n2389, C2 => n2187, ZN => n1525);
   U2058 : OAI222_X1 port map( A1 => n2294, A2 => n2387, B1 => n3158, B2 => 
                           n2388, C1 => n2389, C2 => n2188, ZN => n1524);
   U2059 : OAI222_X1 port map( A1 => n2295, A2 => n2387, B1 => n3146, B2 => 
                           n2388, C1 => n2389, C2 => n2189, ZN => n1523);
   U2060 : OAI222_X1 port map( A1 => n2296, A2 => n2387, B1 => n3134, B2 => 
                           n2388, C1 => n2389, C2 => n2190, ZN => n1522);
   U2061 : OAI222_X1 port map( A1 => n2297, A2 => n2387, B1 => n3122, B2 => 
                           n2388, C1 => n2389, C2 => n2191, ZN => n1521);
   U2062 : OAI222_X1 port map( A1 => n2298, A2 => n2387, B1 => n3112, B2 => 
                           n2388, C1 => n2389, C2 => n2192, ZN => n1520);
   U2063 : INV_X1 port map( A => n2390, ZN => n2389);
   U2064 : AND3_X1 port map( A1 => n2390, A2 => n2300, A3 => n2369, ZN => n2388
                           );
   U2065 : NAND2_X1 port map( A1 => n2199, A2 => n2234, ZN => n2300);
   U2066 : NAND3_X1 port map( A1 => n2235, A2 => n2390, A3 => n2371, ZN => 
                           n2387);
   U2067 : OAI21_X1 port map( B1 => n2219, B2 => n2391, A => n2181, ZN => n2390
                           );
   U2068 : INV_X1 port map( A => n2234, ZN => n2235);
   U2069 : NAND3_X1 port map( A1 => N1662, A2 => n2149, A3 => N1663, ZN => 
                           n2234);
   U2070 : OAI222_X1 port map( A1 => n2290, A2 => n2392, B1 => n2393, B2 => 
                           n1882, C1 => n2394, C2 => n2185, ZN => n1519);
   U2071 : OAI222_X1 port map( A1 => n2292, A2 => n2392, B1 => n2393, B2 => 
                           n1883, C1 => n2394, C2 => n2186, ZN => n1518);
   U2072 : OAI222_X1 port map( A1 => n2293, A2 => n2392, B1 => n2393, B2 => 
                           n1884, C1 => n2394, C2 => n2187, ZN => n1517);
   U2073 : OAI222_X1 port map( A1 => n2294, A2 => n2392, B1 => n2393, B2 => 
                           n1885, C1 => n2394, C2 => n2188, ZN => n1516);
   U2074 : OAI222_X1 port map( A1 => n2295, A2 => n2392, B1 => n2393, B2 => 
                           n1886, C1 => n2394, C2 => n2189, ZN => n1515);
   U2075 : OAI222_X1 port map( A1 => n2296, A2 => n2392, B1 => n2393, B2 => 
                           n1887, C1 => n2394, C2 => n2190, ZN => n1514);
   U2076 : OAI222_X1 port map( A1 => n2297, A2 => n2392, B1 => n2393, B2 => 
                           n1888, C1 => n2394, C2 => n2191, ZN => n1513);
   U2077 : OAI222_X1 port map( A1 => n2298, A2 => n2392, B1 => n2393, B2 => 
                           n1807, C1 => n2394, C2 => n2192, ZN => n1512);
   U2078 : INV_X1 port map( A => n2395, ZN => n2394);
   U2079 : AND3_X1 port map( A1 => n2395, A2 => n2307, A3 => n2369, ZN => n2393
                           );
   U2080 : NAND2_X1 port map( A1 => n2199, A2 => n2241, ZN => n2307);
   U2081 : NAND3_X1 port map( A1 => n2242, A2 => n2395, A3 => n2371, ZN => 
                           n2392);
   U2082 : OAI21_X1 port map( B1 => n2243, B2 => n2377, A => n2181, ZN => n2395
                           );
   U2083 : NAND2_X1 port map( A1 => n2259, A2 => n2396, ZN => n2377);
   U2084 : INV_X1 port map( A => n2219, ZN => n2259);
   U2085 : INV_X1 port map( A => n2241, ZN => n2242);
   U2086 : NAND3_X1 port map( A1 => n2147, A2 => n2149, A3 => N1663, ZN => 
                           n2241);
   U2087 : OAI222_X1 port map( A1 => n2290, A2 => n2397, B1 => n3195, B2 => 
                           n2398, C1 => n2399, C2 => n2185, ZN => n1511);
   U2088 : OAI222_X1 port map( A1 => n2292, A2 => n2397, B1 => n3183, B2 => 
                           n2398, C1 => n2399, C2 => n2186, ZN => n1510);
   U2089 : OAI222_X1 port map( A1 => n2293, A2 => n2397, B1 => n3171, B2 => 
                           n2398, C1 => n2399, C2 => n2187, ZN => n1509);
   U2090 : OAI222_X1 port map( A1 => n2294, A2 => n2397, B1 => n3159, B2 => 
                           n2398, C1 => n2399, C2 => n2188, ZN => n1508);
   U2091 : OAI222_X1 port map( A1 => n2295, A2 => n2397, B1 => n3147, B2 => 
                           n2398, C1 => n2399, C2 => n2189, ZN => n1507);
   U2092 : OAI222_X1 port map( A1 => n2296, A2 => n2397, B1 => n3135, B2 => 
                           n2398, C1 => n2399, C2 => n2190, ZN => n1506);
   U2093 : OAI222_X1 port map( A1 => n2297, A2 => n2397, B1 => n3123, B2 => 
                           n2398, C1 => n2399, C2 => n2191, ZN => n1505);
   U2094 : OAI222_X1 port map( A1 => n2298, A2 => n2397, B1 => n3113, B2 => 
                           n2398, C1 => n2399, C2 => n2192, ZN => n1504);
   U2095 : INV_X1 port map( A => n2400, ZN => n2399);
   U2096 : AND3_X1 port map( A1 => n2400, A2 => n2311, A3 => n2369, ZN => n2398
                           );
   U2097 : NAND2_X1 port map( A1 => n2199, A2 => n2249, ZN => n2311);
   U2098 : NAND3_X1 port map( A1 => n2250, A2 => n2400, A3 => n2371, ZN => 
                           n2397);
   U2099 : OAI21_X1 port map( B1 => n2219, B2 => n2401, A => n2181, ZN => n2400
                           );
   U2100 : INV_X1 port map( A => n2249, ZN => n2250);
   U2101 : NAND3_X1 port map( A1 => n2148, A2 => n2149, A3 => N1662, ZN => 
                           n2249);
   U2102 : OAI222_X1 port map( A1 => n2290, A2 => n2402, B1 => n2185, B2 => 
                           n2403, C1 => n2404, C2 => n1998, ZN => n1503);
   U2103 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(0), ZN => n2290);
   U2104 : OAI222_X1 port map( A1 => n2292, A2 => n2402, B1 => n2186, B2 => 
                           n2403, C1 => n2404, C2 => n1999, ZN => n1502);
   U2105 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(1), ZN => n2292);
   U2106 : OAI222_X1 port map( A1 => n2293, A2 => n2402, B1 => n2187, B2 => 
                           n2403, C1 => n2404, C2 => n2000, ZN => n1501);
   U2107 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(2), ZN => n2293);
   U2108 : OAI222_X1 port map( A1 => n2294, A2 => n2402, B1 => n2188, B2 => 
                           n2403, C1 => n2404, C2 => n2001, ZN => n1500);
   U2109 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(3), ZN => n2294);
   U2110 : OAI222_X1 port map( A1 => n2295, A2 => n2402, B1 => n2189, B2 => 
                           n2403, C1 => n2404, C2 => n2002, ZN => n1499);
   U2111 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(4), ZN => n2295);
   U2112 : OAI222_X1 port map( A1 => n2296, A2 => n2402, B1 => n2190, B2 => 
                           n2403, C1 => n2404, C2 => n2003, ZN => n1498);
   U2113 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(5), ZN => n2296);
   U2114 : OAI222_X1 port map( A1 => n2297, A2 => n2402, B1 => n2191, B2 => 
                           n2403, C1 => n2404, C2 => n2004, ZN => n1497);
   U2115 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(6), ZN => n2297);
   U2116 : OAI222_X1 port map( A1 => n2404, A2 => n1997, B1 => n2192, B2 => 
                           n2403, C1 => n2298, C2 => n2402, ZN => n1496);
   U2117 : NAND3_X1 port map( A1 => n2371, A2 => n2258, A3 => n2406, ZN => 
                           n2402);
   U2118 : INV_X1 port map( A => n2257, ZN => n2258);
   U2119 : NAND2_X1 port map( A1 => n2260, A2 => DATAIN(7), ZN => n2298);
   U2120 : NOR2_X1 port map( A1 => n2132, A2 => n2407, ZN => n2260);
   U2121 : INV_X1 port map( A => n2133, ZN => n2405);
   U2122 : AND3_X1 port map( A1 => n2369, A2 => n2318, A3 => n2406, ZN => n2404
                           );
   U2123 : INV_X1 port map( A => n2403, ZN => n2406);
   U2124 : OAI21_X1 port map( B1 => n2127, B2 => n2201, A => n2202, ZN => n2403
                           );
   U2125 : NAND2_X1 port map( A1 => n2181, A2 => n2219, ZN => n2202);
   U2126 : NAND3_X1 port map( A1 => n2137, A2 => n1266, A3 => n2138, ZN => 
                           n2219);
   U2127 : NAND2_X1 port map( A1 => n3286, A2 => n3283, ZN => n2138);
   U2128 : INV_X1 port map( A => n2408, ZN => n2137);
   U2129 : INV_X1 port map( A => n2181, ZN => n2201);
   U2130 : NAND2_X1 port map( A1 => n2199, A2 => n2257, ZN => n2318);
   U2131 : NAND3_X1 port map( A1 => n2148, A2 => n2149, A3 => n2147, ZN => 
                           n2257);
   U2132 : INV_X1 port map( A => N1662, ZN => n2147);
   U2133 : INV_X1 port map( A => N1664, ZN => n2149);
   U2134 : INV_X1 port map( A => N1663, ZN => n2148);
   U2135 : INV_X1 port map( A => n2410, ZN => n2369);
   U2136 : OAI21_X1 port map( B1 => n2371, B2 => n2132, A => n2320, ZN => n2410
                           );
   U2137 : NAND2_X1 port map( A1 => n2407, A2 => n2199, ZN => n2320);
   U2138 : INV_X1 port map( A => n2132, ZN => n2199);
   U2139 : INV_X1 port map( A => n2180, ZN => n2407);
   U2140 : NOR2_X1 port map( A1 => N1665, A2 => N1666, ZN => n2371);
   U2141 : NAND4_X1 port map( A1 => n2411, A2 => n2412, A3 => n2413, A4 => 
                           n2414, ZN => n1273);
   U2142 : AOI221_X1 port map( B1 => n2128, B2 => n2415, C1 => n2127, C2 => 
                           n3280, A => n2416, ZN => n2414);
   U2143 : OAI222_X1 port map( A1 => n2417, A2 => n2418, B1 => n2419, B2 => 
                           n2420, C1 => n2421, C2 => n2422, ZN => n2416);
   U2144 : AOI221_X1 port map( B1 => n3076, B2 => n2129, C1 => n3192, C2 => 
                           n2423, A => n2424, ZN => n2421);
   U2145 : OAI22_X1 port map( A1 => n3191, A2 => n2115, B1 => n2274, B2 => 
                           n1911, ZN => n2424);
   U2146 : INV_X1 port map( A => n2425, ZN => n2419);
   U2147 : OAI222_X1 port map( A1 => n2274, A2 => n3196, B1 => n2243, B2 => 
                           n3195, C1 => n2228, C2 => n3194, ZN => n2425);
   U2148 : AOI221_X1 port map( B1 => n2426, B2 => n1902, C1 => n2427, C2 => 
                           n1842, A => n2428, ZN => n2417);
   U2149 : OAI22_X1 port map( A1 => n3029, A2 => n2274, B1 => n3274, B2 => 
                           n2339, ZN => n2428);
   U2150 : OAI221_X1 port map( B1 => n2228, B2 => n1800, C1 => n2115, C2 => 
                           n1925, A => n2429, ZN => n2415);
   U2151 : AOI222_X1 port map( A1 => n3084, A2 => n2427, B1 => n3092, B2 => 
                           n2423, C1 => n3217, C2 => n2426, ZN => n2429);
   U2152 : AOI221_X1 port map( B1 => n2365, B2 => n3278, C1 => n2372, C2 => 
                           n3052, A => n2430, ZN => n2413);
   U2153 : OAI222_X1 port map( A1 => n2401, A2 => n1998, B1 => n2382, B2 => 
                           n1823, C1 => n2391, C2 => n1882, ZN => n2430);
   U2154 : AOI221_X1 port map( B1 => n2302, B2 => n3068, C1 => n2313, C2 => 
                           n3060, A => n2431, ZN => n2412);
   U2155 : OAI222_X1 port map( A1 => n2354, A2 => n1808, B1 => n2126, B2 => 
                           n1981, C1 => n2345, C2 => n1831, ZN => n2431);
   U2156 : AOI221_X1 port map( B1 => n2200, B2 => n3218, C1 => n2210, C2 => 
                           n3100, A => n2432, ZN => n2411);
   U2157 : OAI222_X1 port map( A1 => n2287, A2 => n1873, B1 => n2218, B2 => 
                           n1816, C1 => n2280, C2 => n1988, ZN => n2432);
   U2158 : NAND4_X1 port map( A1 => n2433, A2 => n2434, A3 => n2435, A4 => 
                           n2436, ZN => n1272);
   U2159 : AOI221_X1 port map( B1 => n2128, B2 => n2437, C1 => n2127, C2 => 
                           n3272, A => n2438, ZN => n2436);
   U2160 : OAI222_X1 port map( A1 => n2439, A2 => n2418, B1 => n2440, B2 => 
                           n2420, C1 => n2441, C2 => n2422, ZN => n2438);
   U2161 : AOI221_X1 port map( B1 => n3075, B2 => n2129, C1 => n3180, C2 => 
                           n2423, A => n2442, ZN => n2441);
   U2162 : OAI22_X1 port map( A1 => n3179, A2 => n2115, B1 => n2274, B2 => 
                           n1912, ZN => n2442);
   U2163 : INV_X1 port map( A => n2443, ZN => n2440);
   U2164 : OAI222_X1 port map( A1 => n2274, A2 => n3184, B1 => n2243, B2 => 
                           n3183, C1 => n2228, C2 => n3182, ZN => n2443);
   U2165 : AOI221_X1 port map( B1 => n2426, B2 => n1903, C1 => n2427, C2 => 
                           n1843, A => n2444, ZN => n2439);
   U2166 : OAI22_X1 port map( A1 => n3030, A2 => n2274, B1 => n3266, B2 => 
                           n2339, ZN => n2444);
   U2167 : OAI221_X1 port map( B1 => n2228, B2 => n1801, C1 => n2115, C2 => 
                           n1926, A => n2445, ZN => n2437);
   U2168 : AOI222_X1 port map( A1 => n3083, A2 => n2427, B1 => n3091, B2 => 
                           n2423, C1 => n3215, C2 => n2426, ZN => n2445);
   U2169 : AOI221_X1 port map( B1 => n2365, B2 => n3270, C1 => n2372, C2 => 
                           n3051, A => n2446, ZN => n2435);
   U2170 : OAI222_X1 port map( A1 => n2401, A2 => n1999, B1 => n2382, B2 => 
                           n1824, C1 => n2391, C2 => n1883, ZN => n2446);
   U2171 : AOI221_X1 port map( B1 => n2302, B2 => n3067, C1 => n2313, C2 => 
                           n3059, A => n2447, ZN => n2434);
   U2172 : OAI222_X1 port map( A1 => n2354, A2 => n1809, B1 => n2126, B2 => 
                           n1982, C1 => n2345, C2 => n1832, ZN => n2447);
   U2173 : AOI221_X1 port map( B1 => n2200, B2 => n3216, C1 => n2210, C2 => 
                           n3099, A => n2448, ZN => n2433);
   U2174 : OAI222_X1 port map( A1 => n2287, A2 => n1874, B1 => n2218, B2 => 
                           n1817, C1 => n2280, C2 => n1989, ZN => n2448);
   U2175 : NAND4_X1 port map( A1 => n2449, A2 => n2450, A3 => n2451, A4 => 
                           n2452, ZN => n1271);
   U2176 : AOI221_X1 port map( B1 => n2128, B2 => n2453, C1 => n2127, C2 => 
                           n3264, A => n2454, ZN => n2452);
   U2177 : OAI222_X1 port map( A1 => n2455, A2 => n2418, B1 => n2456, B2 => 
                           n2420, C1 => n2457, C2 => n2422, ZN => n2454);
   U2178 : AOI221_X1 port map( B1 => n3074, B2 => n2129, C1 => n3168, C2 => 
                           n2423, A => n2458, ZN => n2457);
   U2179 : OAI22_X1 port map( A1 => n3167, A2 => n2115, B1 => n2274, B2 => 
                           n1913, ZN => n2458);
   U2180 : INV_X1 port map( A => n2459, ZN => n2456);
   U2181 : OAI222_X1 port map( A1 => n2274, A2 => n3172, B1 => n2243, B2 => 
                           n3171, C1 => n2228, C2 => n3170, ZN => n2459);
   U2182 : AOI221_X1 port map( B1 => n2426, B2 => n1904, C1 => n2427, C2 => 
                           n1844, A => n2460, ZN => n2455);
   U2183 : OAI22_X1 port map( A1 => n3031, A2 => n2274, B1 => n3258, B2 => 
                           n2339, ZN => n2460);
   U2184 : OAI221_X1 port map( B1 => n2228, B2 => n1802, C1 => n2115, C2 => 
                           n1927, A => n2461, ZN => n2453);
   U2185 : AOI222_X1 port map( A1 => n3082, A2 => n2427, B1 => n3090, B2 => 
                           n2423, C1 => n3213, C2 => n2426, ZN => n2461);
   U2186 : AOI221_X1 port map( B1 => n2365, B2 => n3262, C1 => n2372, C2 => 
                           n3050, A => n2462, ZN => n2451);
   U2187 : OAI222_X1 port map( A1 => n2401, A2 => n2000, B1 => n2382, B2 => 
                           n1825, C1 => n2391, C2 => n1884, ZN => n2462);
   U2188 : AOI221_X1 port map( B1 => n2302, B2 => n3066, C1 => n2313, C2 => 
                           n3058, A => n2463, ZN => n2450);
   U2189 : OAI222_X1 port map( A1 => n2354, A2 => n1810, B1 => n2126, B2 => 
                           n1983, C1 => n2345, C2 => n1833, ZN => n2463);
   U2190 : AOI221_X1 port map( B1 => n2200, B2 => n3214, C1 => n2210, C2 => 
                           n3098, A => n2464, ZN => n2449);
   U2191 : OAI222_X1 port map( A1 => n2287, A2 => n1875, B1 => n2218, B2 => 
                           n1818, C1 => n2280, C2 => n1990, ZN => n2464);
   U2192 : NAND4_X1 port map( A1 => n2465, A2 => n2466, A3 => n2467, A4 => 
                           n2468, ZN => n1270);
   U2193 : AOI221_X1 port map( B1 => n2128, B2 => n2469, C1 => n2127, C2 => 
                           n3256, A => n2470, ZN => n2468);
   U2194 : OAI222_X1 port map( A1 => n2471, A2 => n2418, B1 => n2472, B2 => 
                           n2420, C1 => n2473, C2 => n2422, ZN => n2470);
   U2195 : AOI221_X1 port map( B1 => n3073, B2 => n2129, C1 => n3156, C2 => 
                           n2423, A => n2474, ZN => n2473);
   U2196 : OAI22_X1 port map( A1 => n3155, A2 => n2115, B1 => n2274, B2 => 
                           n1914, ZN => n2474);
   U2197 : INV_X1 port map( A => n2475, ZN => n2472);
   U2198 : OAI222_X1 port map( A1 => n2274, A2 => n3160, B1 => n2243, B2 => 
                           n3159, C1 => n2228, C2 => n3158, ZN => n2475);
   U2199 : AOI221_X1 port map( B1 => n2426, B2 => n1905, C1 => n2427, C2 => 
                           n1845, A => n2476, ZN => n2471);
   U2200 : OAI22_X1 port map( A1 => n3032, A2 => n2274, B1 => n3250, B2 => 
                           n2339, ZN => n2476);
   U2201 : OAI221_X1 port map( B1 => n2228, B2 => n1803, C1 => n2115, C2 => 
                           n1928, A => n2477, ZN => n2469);
   U2202 : AOI222_X1 port map( A1 => n3081, A2 => n2427, B1 => n3089, B2 => 
                           n2423, C1 => n3211, C2 => n2426, ZN => n2477);
   U2203 : AOI221_X1 port map( B1 => n2365, B2 => n3254, C1 => n2372, C2 => 
                           n3049, A => n2478, ZN => n2467);
   U2204 : OAI222_X1 port map( A1 => n2401, A2 => n2001, B1 => n2382, B2 => 
                           n1826, C1 => n2391, C2 => n1885, ZN => n2478);
   U2205 : AOI221_X1 port map( B1 => n2302, B2 => n3065, C1 => n2313, C2 => 
                           n3057, A => n2479, ZN => n2466);
   U2206 : OAI222_X1 port map( A1 => n2354, A2 => n1811, B1 => n2126, B2 => 
                           n1984, C1 => n2345, C2 => n1834, ZN => n2479);
   U2207 : AOI221_X1 port map( B1 => n2200, B2 => n3212, C1 => n2210, C2 => 
                           n3097, A => n2480, ZN => n2465);
   U2208 : OAI222_X1 port map( A1 => n2287, A2 => n1876, B1 => n2218, B2 => 
                           n1819, C1 => n2280, C2 => n1991, ZN => n2480);
   U2209 : NAND4_X1 port map( A1 => n2481, A2 => n2482, A3 => n2483, A4 => 
                           n2484, ZN => n1269);
   U2210 : AOI221_X1 port map( B1 => n2128, B2 => n2485, C1 => n2127, C2 => 
                           n3248, A => n2486, ZN => n2484);
   U2211 : OAI222_X1 port map( A1 => n2487, A2 => n2418, B1 => n2488, B2 => 
                           n2420, C1 => n2489, C2 => n2422, ZN => n2486);
   U2212 : AOI221_X1 port map( B1 => n3072, B2 => n2129, C1 => n3144, C2 => 
                           n2423, A => n2490, ZN => n2489);
   U2213 : OAI22_X1 port map( A1 => n3143, A2 => n2115, B1 => n2274, B2 => 
                           n1915, ZN => n2490);
   U2214 : INV_X1 port map( A => n2491, ZN => n2488);
   U2215 : OAI222_X1 port map( A1 => n2274, A2 => n3148, B1 => n2243, B2 => 
                           n3147, C1 => n2228, C2 => n3146, ZN => n2491);
   U2216 : AOI221_X1 port map( B1 => n2426, B2 => n1906, C1 => n2427, C2 => 
                           n1846, A => n2492, ZN => n2487);
   U2217 : OAI22_X1 port map( A1 => n3033, A2 => n2274, B1 => n3242, B2 => 
                           n2339, ZN => n2492);
   U2218 : OAI221_X1 port map( B1 => n2228, B2 => n1804, C1 => n2115, C2 => 
                           n1929, A => n2493, ZN => n2485);
   U2219 : AOI222_X1 port map( A1 => n3080, A2 => n2427, B1 => n3088, B2 => 
                           n2423, C1 => n3209, C2 => n2426, ZN => n2493);
   U2220 : AOI221_X1 port map( B1 => n2365, B2 => n3246, C1 => n2372, C2 => 
                           n3048, A => n2494, ZN => n2483);
   U2221 : OAI222_X1 port map( A1 => n2401, A2 => n2002, B1 => n2382, B2 => 
                           n1827, C1 => n2391, C2 => n1886, ZN => n2494);
   U2222 : AOI221_X1 port map( B1 => n2302, B2 => n3064, C1 => n2313, C2 => 
                           n3056, A => n2495, ZN => n2482);
   U2223 : OAI222_X1 port map( A1 => n2354, A2 => n1812, B1 => n2126, B2 => 
                           n1985, C1 => n2345, C2 => n1835, ZN => n2495);
   U2224 : AOI221_X1 port map( B1 => n2200, B2 => n3210, C1 => n2210, C2 => 
                           n3096, A => n2496, ZN => n2481);
   U2225 : OAI222_X1 port map( A1 => n2287, A2 => n1877, B1 => n2218, B2 => 
                           n1820, C1 => n2280, C2 => n1992, ZN => n2496);
   U2226 : NAND4_X1 port map( A1 => n2497, A2 => n2498, A3 => n2499, A4 => 
                           n2500, ZN => n1268);
   U2227 : AOI221_X1 port map( B1 => n2128, B2 => n2501, C1 => n2127, C2 => 
                           n3240, A => n2502, ZN => n2500);
   U2228 : OAI222_X1 port map( A1 => n2503, A2 => n2418, B1 => n2504, B2 => 
                           n2420, C1 => n2505, C2 => n2422, ZN => n2502);
   U2229 : AOI221_X1 port map( B1 => n3071, B2 => n2129, C1 => n3132, C2 => 
                           n2423, A => n2506, ZN => n2505);
   U2230 : OAI22_X1 port map( A1 => n3131, A2 => n2115, B1 => n2274, B2 => 
                           n1916, ZN => n2506);
   U2231 : INV_X1 port map( A => n2507, ZN => n2504);
   U2232 : OAI222_X1 port map( A1 => n2274, A2 => n3136, B1 => n2243, B2 => 
                           n3135, C1 => n2228, C2 => n3134, ZN => n2507);
   U2233 : AOI221_X1 port map( B1 => n2426, B2 => n1892, C1 => n2427, C2 => 
                           n1847, A => n2508, ZN => n2503);
   U2234 : OAI22_X1 port map( A1 => n3034, A2 => n2274, B1 => n3234, B2 => 
                           n2339, ZN => n2508);
   U2235 : OAI221_X1 port map( B1 => n2228, B2 => n1805, C1 => n2115, C2 => 
                           n1930, A => n2509, ZN => n2501);
   U2236 : AOI222_X1 port map( A1 => n3079, A2 => n2427, B1 => n3087, B2 => 
                           n2423, C1 => n3207, C2 => n2426, ZN => n2509);
   U2237 : AOI221_X1 port map( B1 => n2365, B2 => n3238, C1 => n2372, C2 => 
                           n3047, A => n2510, ZN => n2499);
   U2238 : OAI222_X1 port map( A1 => n2401, A2 => n2003, B1 => n2382, B2 => 
                           n1828, C1 => n2391, C2 => n1887, ZN => n2510);
   U2239 : AOI221_X1 port map( B1 => n2302, B2 => n3063, C1 => n2313, C2 => 
                           n3055, A => n2511, ZN => n2498);
   U2240 : OAI222_X1 port map( A1 => n2354, A2 => n1813, B1 => n2126, B2 => 
                           n1986, C1 => n2345, C2 => n1836, ZN => n2511);
   U2241 : AOI221_X1 port map( B1 => n2200, B2 => n3208, C1 => n2210, C2 => 
                           n3095, A => n2512, ZN => n2497);
   U2242 : OAI222_X1 port map( A1 => n2287, A2 => n1878, B1 => n2218, B2 => 
                           n1821, C1 => n2280, C2 => n1993, ZN => n2512);
   U2243 : NAND4_X1 port map( A1 => n2513, A2 => n2514, A3 => n2515, A4 => 
                           n2516, ZN => n1267);
   U2244 : AOI221_X1 port map( B1 => n2128, B2 => n2517, C1 => n2127, C2 => 
                           n3232, A => n2518, ZN => n2516);
   U2245 : OAI222_X1 port map( A1 => n2519, A2 => n2418, B1 => n2520, B2 => 
                           n2420, C1 => n2521, C2 => n2422, ZN => n2518);
   U2246 : AOI221_X1 port map( B1 => n3070, B2 => n2129, C1 => n3120, C2 => 
                           n2423, A => n2522, ZN => n2521);
   U2247 : OAI22_X1 port map( A1 => n3119, A2 => n2115, B1 => n2274, B2 => 
                           n1917, ZN => n2522);
   U2248 : INV_X1 port map( A => n2523, ZN => n2520);
   U2249 : OAI222_X1 port map( A1 => n2274, A2 => n3124, B1 => n2243, B2 => 
                           n3123, C1 => n2228, C2 => n3122, ZN => n2523);
   U2250 : AOI221_X1 port map( B1 => n2426, B2 => n1893, C1 => n2427, C2 => 
                           n1841, A => n2524, ZN => n2519);
   U2251 : OAI22_X1 port map( A1 => n3035, A2 => n2274, B1 => n3226, B2 => 
                           n2339, ZN => n2524);
   U2252 : OAI221_X1 port map( B1 => n2228, B2 => n1806, C1 => n2115, C2 => 
                           n1931, A => n2525, ZN => n2517);
   U2253 : AOI222_X1 port map( A1 => n3078, A2 => n2427, B1 => n3086, B2 => 
                           n2423, C1 => n3205, C2 => n2426, ZN => n2525);
   U2254 : AOI221_X1 port map( B1 => n2365, B2 => n3230, C1 => n2372, C2 => 
                           n3046, A => n2526, ZN => n2515);
   U2255 : OAI222_X1 port map( A1 => n2401, A2 => n2004, B1 => n2382, B2 => 
                           n1829, C1 => n2391, C2 => n1888, ZN => n2526);
   U2256 : AOI221_X1 port map( B1 => n2302, B2 => n3062, C1 => n2313, C2 => 
                           n3054, A => n2527, ZN => n2514);
   U2257 : OAI222_X1 port map( A1 => n2354, A2 => n1814, B1 => n2126, B2 => 
                           n1987, C1 => n2345, C2 => n1837, ZN => n2527);
   U2258 : AOI221_X1 port map( B1 => n2200, B2 => n3206, C1 => n2210, C2 => 
                           n3094, A => n2528, ZN => n2513);
   U2259 : OAI222_X1 port map( A1 => n2287, A2 => n1879, B1 => n2218, B2 => 
                           n1822, C1 => n2280, C2 => n1994, ZN => n2528);
   U2260 : NAND4_X1 port map( A1 => n2529, A2 => n2530, A3 => n2531, A4 => 
                           n2532, ZN => n1265);
   U2261 : AOI221_X1 port map( B1 => n2128, B2 => n2533, C1 => n2127, C2 => 
                           n3224, A => n2534, ZN => n2532);
   U2262 : OAI222_X1 port map( A1 => n2535, A2 => n2418, B1 => n2536, B2 => 
                           n2420, C1 => n2537, C2 => n2422, ZN => n2534);
   U2263 : AOI221_X1 port map( B1 => n3069, B2 => n2129, C1 => n3110, C2 => 
                           n2423, A => n2538, ZN => n2537);
   U2264 : OAI22_X1 port map( A1 => n3109, A2 => n2115, B1 => n2274, B2 => 
                           n1871, ZN => n2538);
   U2265 : INV_X1 port map( A => n2539, ZN => n2536);
   U2266 : OAI222_X1 port map( A1 => n2274, A2 => n3114, B1 => n2243, B2 => 
                           n3113, C1 => n2228, C2 => n3112, ZN => n2539);
   U2267 : AOI221_X1 port map( B1 => n2426, B2 => n2005, C1 => n2427, C2 => 
                           n1840, A => n2540, ZN => n2535);
   U2268 : OAI22_X1 port map( A1 => n3036, A2 => n2274, B1 => n3220, B2 => 
                           n2339, ZN => n2540);
   U2269 : NOR2_X1 port map( A1 => n2420, A2 => n2115, ZN => n2127);
   U2270 : OAI221_X1 port map( B1 => n2228, B2 => n1890, C1 => n2115, C2 => 
                           n1839, A => n2541, ZN => n2533);
   U2271 : AOI222_X1 port map( A1 => n3077, A2 => n2427, B1 => n3085, B2 => 
                           n2423, C1 => n3203, C2 => n2426, ZN => n2541);
   U2272 : INV_X1 port map( A => n2542, ZN => n2228);
   U2273 : AOI221_X1 port map( B1 => n2365, B2 => n3223, C1 => n2372, C2 => 
                           n3045, A => n2543, ZN => n2531);
   U2274 : OAI222_X1 port map( A1 => n2401, A2 => n1997, B1 => n2382, B2 => 
                           n1881, C1 => n2391, C2 => n1807, ZN => n2543);
   U2275 : NAND2_X1 port map( A1 => n2396, A2 => n2426, ZN => n2391);
   U2276 : INV_X1 port map( A => n2113, ZN => n2426);
   U2277 : NAND2_X1 port map( A1 => n2544, A2 => n2396, ZN => n2382);
   U2278 : NAND2_X1 port map( A1 => n2427, A2 => n2396, ZN => n2401);
   U2279 : INV_X1 port map( A => n2420, ZN => n2396);
   U2280 : INV_X1 port map( A => n2251, ZN => n2427);
   U2281 : NOR2_X1 port map( A1 => n2420, A2 => n2120, ZN => n2372);
   U2282 : NAND2_X1 port map( A1 => n1491, A2 => n1492, ZN => n2420);
   U2283 : NOR2_X1 port map( A1 => n2418, A2 => n2115, ZN => n2365);
   U2284 : AOI221_X1 port map( B1 => n2302, B2 => n3061, C1 => n2313, C2 => 
                           n3053, A => n2545, ZN => n2530);
   U2285 : OAI222_X1 port map( A1 => n2354, A2 => n1891, B1 => n2126, B2 => 
                           n1799, C1 => n2345, C2 => n1838, ZN => n2545);
   U2286 : NAND2_X1 port map( A1 => n2542, A2 => n2359, ZN => n2345);
   U2287 : NAND2_X1 port map( A1 => n2359, A2 => n2129, ZN => n2126);
   U2288 : INV_X1 port map( A => n2120, ZN => n2129);
   U2289 : NAND2_X1 port map( A1 => n2423, A2 => n2359, ZN => n2354);
   U2290 : INV_X1 port map( A => n2418, ZN => n2359);
   U2291 : NAND2_X1 port map( A1 => n1491, A2 => n1934, ZN => n2418);
   U2292 : INV_X1 port map( A => n2243, ZN => n2423);
   U2293 : NAND3_X1 port map( A1 => n1495, A2 => n1830, A3 => n1493, ZN => 
                           n2243);
   U2294 : NOR2_X1 port map( A1 => n2422, A2 => n2251, ZN => n2313);
   U2295 : NAND3_X1 port map( A1 => n1494, A2 => n1798, A3 => n1493, ZN => 
                           n2251);
   U2296 : NOR2_X1 port map( A1 => n2422, A2 => n2113, ZN => n2302);
   U2297 : NAND3_X1 port map( A1 => n1830, A2 => n1798, A3 => n1493, ZN => 
                           n2113);
   U2298 : INV_X1 port map( A => n2125, ZN => n2422);
   U2299 : AOI221_X1 port map( B1 => n2200, B2 => n3204, C1 => n2210, C2 => 
                           n3093, A => n2546, ZN => n2529);
   U2300 : OAI222_X1 port map( A1 => n2287, A2 => n1815, B1 => n2218, B2 => 
                           n1880, C1 => n2280, C2 => n1995, ZN => n2546);
   U2301 : NAND2_X1 port map( A1 => n2125, A2 => n2544, ZN => n2280);
   U2302 : NAND2_X1 port map( A1 => n2544, A2 => n2128, ZN => n2218);
   U2303 : INV_X1 port map( A => n2339, ZN => n2544);
   U2304 : NAND3_X1 port map( A1 => n1889, A2 => n1798, A3 => n1494, ZN => 
                           n2339);
   U2305 : NAND2_X1 port map( A1 => n2125, A2 => n2542, ZN => n2287);
   U2306 : NOR2_X1 port map( A1 => n2111, A2 => n1493, ZN => n2542);
   U2307 : NOR2_X1 port map( A1 => n1934, A2 => n1491, ZN => n2125);
   U2308 : NOR2_X1 port map( A1 => n2274, A2 => n2547, ZN => n2210);
   U2309 : NOR2_X1 port map( A1 => n2547, A2 => n2120, ZN => n2200);
   U2310 : NAND3_X1 port map( A1 => n1830, A2 => n1798, A3 => n1889, ZN => 
                           n2120);
   U2311 : INV_X1 port map( A => n2128, ZN => n2547);
   U2312 : NOR2_X1 port map( A1 => n1491, A2 => n1492, ZN => n2128);
   U2313 : NAND2_X1 port map( A1 => n2548, A2 => n2549, ZN => n1264);
   U2314 : NOR4_X1 port map( A1 => n2550, A2 => n2551, A3 => n2552, A4 => n2553
                           , ZN => n2549);
   U2315 : AOI21_X1 port map( B1 => n2554, B2 => n2555, A => n2556, ZN => n2553
                           );
   U2316 : AOI221_X1 port map( B1 => n2557, B2 => n1842, C1 => n2558, C2 => 
                           n3198, A => n2559, ZN => n2555);
   U2317 : OAI22_X1 port map( A1 => n3195, A2 => n2560, B1 => n1808, B2 => 
                           n2561, ZN => n2559);
   U2318 : AOI221_X1 port map( B1 => n2562, B2 => n3060, C1 => n2563, C2 => 
                           n3192, A => n2564, ZN => n2554);
   U2319 : OAI22_X1 port map( A1 => n1966, A2 => n2565, B1 => n1850, B2 => 
                           n2566, ZN => n2564);
   U2320 : AOI21_X1 port map( B1 => n2567, B2 => n2568, A => n2569, ZN => n2552
                           );
   U2321 : AOI221_X1 port map( B1 => n2557, B2 => n1938, C1 => n2558, C2 => 
                           n3197, A => n2570, ZN => n2568);
   U2322 : OAI22_X1 port map( A1 => n3196, A2 => n2560, B1 => n3029, B2 => 
                           n2561, ZN => n2570);
   U2323 : AOI221_X1 port map( B1 => n2562, B2 => n3202, C1 => n2563, C2 => 
                           n3193, A => n2571, ZN => n2567);
   U2324 : OAI22_X1 port map( A1 => n1816, A2 => n2565, B1 => n1851, B2 => 
                           n2566, ZN => n2571);
   U2325 : AOI21_X1 port map( B1 => n2572, B2 => n2573, A => n2574, ZN => n2551
                           );
   U2326 : AOI221_X1 port map( B1 => n2557, B2 => n3200, C1 => n2558, C2 => 
                           n3052, A => n2575, ZN => n2573);
   U2327 : OAI22_X1 port map( A1 => n1894, A2 => n2560, B1 => n3191, B2 => 
                           n2561, ZN => n2575);
   U2328 : AOI221_X1 port map( B1 => n2562, B2 => n3076, C1 => n2563, C2 => 
                           n3279, A => n2576, ZN => n2572);
   U2329 : OAI22_X1 port map( A1 => n1952, A2 => n2565, B1 => n1864, B2 => 
                           n2566, ZN => n2576);
   U2330 : AOI21_X1 port map( B1 => n2577, B2 => n2578, A => n2579, ZN => n2550
                           );
   U2331 : AOI221_X1 port map( B1 => n2557, B2 => n1902, C1 => n2558, C2 => 
                           n3199, A => n2580, ZN => n2578);
   U2332 : OAI22_X1 port map( A1 => n3194, A2 => n2560, B1 => n1831, B2 => 
                           n2561, ZN => n2580);
   U2333 : AOI221_X1 port map( B1 => n2562, B2 => n3068, C1 => n2563, C2 => 
                           n3277, A => n2581, ZN => n2577);
   U2334 : OAI22_X1 port map( A1 => n1953, A2 => n2565, B1 => n1800, B2 => 
                           n2566, ZN => n2581);
   U2335 : AOI221_X1 port map( B1 => n2582, B2 => n1951, C1 => n2583, C2 => 
                           n3108, A => n2584, ZN => n2548);
   U2336 : OAI22_X1 port map( A1 => n3037, A2 => n2585, B1 => n1918, B2 => 
                           n2586, ZN => n2584);
   U2337 : NAND2_X1 port map( A1 => n2587, A2 => n2588, ZN => n1263);
   U2338 : NOR4_X1 port map( A1 => n2589, A2 => n2590, A3 => n2591, A4 => n2592
                           , ZN => n2588);
   U2339 : AOI21_X1 port map( B1 => n2593, B2 => n2594, A => n2556, ZN => n2592
                           );
   U2340 : AOI221_X1 port map( B1 => n2557, B2 => n1843, C1 => n2558, C2 => 
                           n3186, A => n2595, ZN => n2594);
   U2341 : OAI22_X1 port map( A1 => n3183, A2 => n2560, B1 => n1809, B2 => 
                           n2561, ZN => n2595);
   U2342 : AOI221_X1 port map( B1 => n2562, B2 => n3059, C1 => n2563, C2 => 
                           n3180, A => n2596, ZN => n2593);
   U2343 : OAI22_X1 port map( A1 => n1967, A2 => n2565, B1 => n1852, B2 => 
                           n2566, ZN => n2596);
   U2344 : AOI21_X1 port map( B1 => n2597, B2 => n2598, A => n2569, ZN => n2591
                           );
   U2345 : AOI221_X1 port map( B1 => n2557, B2 => n1939, C1 => n2558, C2 => 
                           n3185, A => n2599, ZN => n2598);
   U2346 : OAI22_X1 port map( A1 => n3184, A2 => n2560, B1 => n3030, B2 => 
                           n2561, ZN => n2599);
   U2347 : AOI221_X1 port map( B1 => n2562, B2 => n3190, C1 => n2563, C2 => 
                           n3181, A => n2600, ZN => n2597);
   U2348 : OAI22_X1 port map( A1 => n1817, A2 => n2565, B1 => n1853, B2 => 
                           n2566, ZN => n2600);
   U2349 : AOI21_X1 port map( B1 => n2601, B2 => n2602, A => n2574, ZN => n2590
                           );
   U2350 : AOI221_X1 port map( B1 => n2557, B2 => n3188, C1 => n2558, C2 => 
                           n3051, A => n2603, ZN => n2602);
   U2351 : OAI22_X1 port map( A1 => n1895, A2 => n2560, B1 => n3179, B2 => 
                           n2561, ZN => n2603);
   U2352 : AOI221_X1 port map( B1 => n2562, B2 => n3075, C1 => n2563, C2 => 
                           n3271, A => n2604, ZN => n2601);
   U2353 : OAI22_X1 port map( A1 => n1954, A2 => n2565, B1 => n1865, B2 => 
                           n2566, ZN => n2604);
   U2354 : AOI21_X1 port map( B1 => n2605, B2 => n2606, A => n2579, ZN => n2589
                           );
   U2355 : AOI221_X1 port map( B1 => n2557, B2 => n1903, C1 => n2558, C2 => 
                           n3187, A => n2607, ZN => n2606);
   U2356 : OAI22_X1 port map( A1 => n3182, A2 => n2560, B1 => n1832, B2 => 
                           n2561, ZN => n2607);
   U2357 : AOI221_X1 port map( B1 => n2562, B2 => n3067, C1 => n2563, C2 => 
                           n3269, A => n2608, ZN => n2605);
   U2358 : OAI22_X1 port map( A1 => n1955, A2 => n2565, B1 => n1801, B2 => 
                           n2566, ZN => n2608);
   U2359 : OAI22_X1 port map( A1 => n3038, A2 => n2585, B1 => n1919, B2 => 
                           n2586, ZN => n2609);
   U2360 : NAND2_X1 port map( A1 => n2610, A2 => n2611, ZN => n1262);
   U2361 : NOR4_X1 port map( A1 => n2612, A2 => n2613, A3 => n2614, A4 => n2615
                           , ZN => n2611);
   U2362 : AOI21_X1 port map( B1 => n2616, B2 => n2617, A => n2556, ZN => n2615
                           );
   U2363 : AOI221_X1 port map( B1 => n2557, B2 => n1844, C1 => n2558, C2 => 
                           n3174, A => n2618, ZN => n2617);
   U2364 : OAI22_X1 port map( A1 => n3171, A2 => n2560, B1 => n1810, B2 => 
                           n2561, ZN => n2618);
   U2365 : AOI221_X1 port map( B1 => n2562, B2 => n3058, C1 => n2563, C2 => 
                           n3168, A => n2619, ZN => n2616);
   U2366 : OAI22_X1 port map( A1 => n1968, A2 => n2565, B1 => n1854, B2 => 
                           n2566, ZN => n2619);
   U2367 : AOI21_X1 port map( B1 => n2620, B2 => n2621, A => n2569, ZN => n2614
                           );
   U2368 : AOI221_X1 port map( B1 => n2557, B2 => n1940, C1 => n2558, C2 => 
                           n3173, A => n2622, ZN => n2621);
   U2369 : OAI22_X1 port map( A1 => n3172, A2 => n2560, B1 => n3031, B2 => 
                           n2561, ZN => n2622);
   U2370 : AOI221_X1 port map( B1 => n2562, B2 => n3178, C1 => n2563, C2 => 
                           n3169, A => n2623, ZN => n2620);
   U2371 : OAI22_X1 port map( A1 => n1818, A2 => n2565, B1 => n1855, B2 => 
                           n2566, ZN => n2623);
   U2372 : AOI21_X1 port map( B1 => n2624, B2 => n2625, A => n2574, ZN => n2613
                           );
   U2373 : AOI221_X1 port map( B1 => n2557, B2 => n3176, C1 => n2558, C2 => 
                           n3050, A => n2626, ZN => n2625);
   U2374 : OAI22_X1 port map( A1 => n1896, A2 => n2560, B1 => n3167, B2 => 
                           n2561, ZN => n2626);
   U2375 : AOI221_X1 port map( B1 => n2562, B2 => n3074, C1 => n2563, C2 => 
                           n3263, A => n2627, ZN => n2624);
   U2376 : OAI22_X1 port map( A1 => n1956, A2 => n2565, B1 => n1866, B2 => 
                           n2566, ZN => n2627);
   U2377 : AOI21_X1 port map( B1 => n2628, B2 => n2629, A => n2579, ZN => n2612
                           );
   U2378 : AOI221_X1 port map( B1 => n2557, B2 => n1904, C1 => n2558, C2 => 
                           n3175, A => n2630, ZN => n2629);
   U2379 : OAI22_X1 port map( A1 => n3170, A2 => n2560, B1 => n1833, B2 => 
                           n2561, ZN => n2630);
   U2380 : AOI221_X1 port map( B1 => n2562, B2 => n3066, C1 => n2563, C2 => 
                           n3261, A => n2631, ZN => n2628);
   U2381 : OAI22_X1 port map( A1 => n1957, A2 => n2565, B1 => n1802, B2 => 
                           n2566, ZN => n2631);
   U2382 : OAI22_X1 port map( A1 => n3039, A2 => n2585, B1 => n1920, B2 => 
                           n2586, ZN => n2632);
   U2383 : NAND2_X1 port map( A1 => n2633, A2 => n2634, ZN => n1261);
   U2384 : NOR4_X1 port map( A1 => n2635, A2 => n2636, A3 => n2637, A4 => n2638
                           , ZN => n2634);
   U2385 : AOI21_X1 port map( B1 => n2639, B2 => n2640, A => n2556, ZN => n2638
                           );
   U2386 : AOI221_X1 port map( B1 => n2557, B2 => n1845, C1 => n2558, C2 => 
                           n3162, A => n2641, ZN => n2640);
   U2387 : OAI22_X1 port map( A1 => n3159, A2 => n2560, B1 => n1811, B2 => 
                           n2561, ZN => n2641);
   U2388 : AOI221_X1 port map( B1 => n2562, B2 => n3057, C1 => n2563, C2 => 
                           n3156, A => n2642, ZN => n2639);
   U2389 : OAI22_X1 port map( A1 => n1969, A2 => n2565, B1 => n1856, B2 => 
                           n2566, ZN => n2642);
   U2390 : AOI21_X1 port map( B1 => n2643, B2 => n2644, A => n2569, ZN => n2637
                           );
   U2391 : AOI221_X1 port map( B1 => n2557, B2 => n1941, C1 => n2558, C2 => 
                           n3161, A => n2645, ZN => n2644);
   U2392 : OAI22_X1 port map( A1 => n3160, A2 => n2560, B1 => n3032, B2 => 
                           n2561, ZN => n2645);
   U2393 : AOI221_X1 port map( B1 => n2562, B2 => n3166, C1 => n2563, C2 => 
                           n3157, A => n2646, ZN => n2643);
   U2394 : OAI22_X1 port map( A1 => n1819, A2 => n2565, B1 => n1857, B2 => 
                           n2566, ZN => n2646);
   U2395 : AOI21_X1 port map( B1 => n2647, B2 => n2648, A => n2574, ZN => n2636
                           );
   U2396 : AOI221_X1 port map( B1 => n2557, B2 => n3164, C1 => n2558, C2 => 
                           n3049, A => n2649, ZN => n2648);
   U2397 : OAI22_X1 port map( A1 => n1897, A2 => n2560, B1 => n3155, B2 => 
                           n2561, ZN => n2649);
   U2398 : AOI221_X1 port map( B1 => n2562, B2 => n3073, C1 => n2563, C2 => 
                           n3255, A => n2650, ZN => n2647);
   U2399 : OAI22_X1 port map( A1 => n1958, A2 => n2565, B1 => n1867, B2 => 
                           n2566, ZN => n2650);
   U2400 : AOI21_X1 port map( B1 => n2651, B2 => n2652, A => n2579, ZN => n2635
                           );
   U2401 : AOI221_X1 port map( B1 => n2557, B2 => n1905, C1 => n2558, C2 => 
                           n3163, A => n2653, ZN => n2652);
   U2402 : OAI22_X1 port map( A1 => n3158, A2 => n2560, B1 => n1834, B2 => 
                           n2561, ZN => n2653);
   U2403 : AOI221_X1 port map( B1 => n2562, B2 => n3065, C1 => n2563, C2 => 
                           n3253, A => n2654, ZN => n2651);
   U2404 : OAI22_X1 port map( A1 => n1959, A2 => n2565, B1 => n1803, B2 => 
                           n2566, ZN => n2654);
   U2405 : OAI22_X1 port map( A1 => n3040, A2 => n2585, B1 => n1921, B2 => 
                           n2586, ZN => n2655);
   U2406 : NAND2_X1 port map( A1 => n2656, A2 => n2657, ZN => n1260);
   U2407 : NOR4_X1 port map( A1 => n2658, A2 => n2659, A3 => n2660, A4 => n2661
                           , ZN => n2657);
   U2408 : AOI21_X1 port map( B1 => n2662, B2 => n2663, A => n2556, ZN => n2661
                           );
   U2409 : AOI221_X1 port map( B1 => n2557, B2 => n1846, C1 => n2558, C2 => 
                           n3150, A => n2664, ZN => n2663);
   U2410 : OAI22_X1 port map( A1 => n3147, A2 => n2560, B1 => n1812, B2 => 
                           n2561, ZN => n2664);
   U2411 : AOI221_X1 port map( B1 => n2562, B2 => n3056, C1 => n2563, C2 => 
                           n3144, A => n2665, ZN => n2662);
   U2412 : OAI22_X1 port map( A1 => n1970, A2 => n2565, B1 => n1858, B2 => 
                           n2566, ZN => n2665);
   U2413 : AOI21_X1 port map( B1 => n2666, B2 => n2667, A => n2569, ZN => n2660
                           );
   U2414 : AOI221_X1 port map( B1 => n2557, B2 => n1942, C1 => n2558, C2 => 
                           n3149, A => n2668, ZN => n2667);
   U2415 : OAI22_X1 port map( A1 => n3148, A2 => n2560, B1 => n3033, B2 => 
                           n2561, ZN => n2668);
   U2416 : AOI221_X1 port map( B1 => n2562, B2 => n3154, C1 => n2563, C2 => 
                           n3145, A => n2669, ZN => n2666);
   U2417 : OAI22_X1 port map( A1 => n1820, A2 => n2565, B1 => n1859, B2 => 
                           n2566, ZN => n2669);
   U2418 : AOI21_X1 port map( B1 => n2670, B2 => n2671, A => n2574, ZN => n2659
                           );
   U2419 : AOI221_X1 port map( B1 => n2557, B2 => n3152, C1 => n2558, C2 => 
                           n3048, A => n2672, ZN => n2671);
   U2420 : OAI22_X1 port map( A1 => n1898, A2 => n2560, B1 => n3143, B2 => 
                           n2561, ZN => n2672);
   U2421 : AOI221_X1 port map( B1 => n2562, B2 => n3072, C1 => n2563, C2 => 
                           n3247, A => n2673, ZN => n2670);
   U2422 : OAI22_X1 port map( A1 => n1960, A2 => n2565, B1 => n1868, B2 => 
                           n2566, ZN => n2673);
   U2423 : AOI21_X1 port map( B1 => n2674, B2 => n2675, A => n2579, ZN => n2658
                           );
   U2424 : AOI221_X1 port map( B1 => n2557, B2 => n1906, C1 => n2558, C2 => 
                           n3151, A => n2676, ZN => n2675);
   U2425 : OAI22_X1 port map( A1 => n3146, A2 => n2560, B1 => n1835, B2 => 
                           n2561, ZN => n2676);
   U2426 : AOI221_X1 port map( B1 => n2562, B2 => n3064, C1 => n2563, C2 => 
                           n3245, A => n2677, ZN => n2674);
   U2427 : OAI22_X1 port map( A1 => n1961, A2 => n2565, B1 => n1804, B2 => 
                           n2566, ZN => n2677);
   U2428 : OAI22_X1 port map( A1 => n3041, A2 => n2585, B1 => n1922, B2 => 
                           n2586, ZN => n2678);
   U2429 : NAND2_X1 port map( A1 => n2679, A2 => n2680, ZN => n1259);
   U2430 : NOR4_X1 port map( A1 => n2681, A2 => n2682, A3 => n2683, A4 => n2684
                           , ZN => n2680);
   U2431 : AOI21_X1 port map( B1 => n2685, B2 => n2686, A => n2556, ZN => n2684
                           );
   U2432 : AOI221_X1 port map( B1 => n2557, B2 => n1847, C1 => n2558, C2 => 
                           n3138, A => n2687, ZN => n2686);
   U2433 : OAI22_X1 port map( A1 => n3135, A2 => n2560, B1 => n1813, B2 => 
                           n2561, ZN => n2687);
   U2434 : AOI221_X1 port map( B1 => n2562, B2 => n3055, C1 => n2563, C2 => 
                           n3132, A => n2688, ZN => n2685);
   U2435 : OAI22_X1 port map( A1 => n1971, A2 => n2565, B1 => n1860, B2 => 
                           n2566, ZN => n2688);
   U2436 : AOI21_X1 port map( B1 => n2689, B2 => n2690, A => n2569, ZN => n2683
                           );
   U2437 : AOI221_X1 port map( B1 => n2557, B2 => n1943, C1 => n2558, C2 => 
                           n3137, A => n2691, ZN => n2690);
   U2438 : OAI22_X1 port map( A1 => n3136, A2 => n2560, B1 => n3034, B2 => 
                           n2561, ZN => n2691);
   U2439 : AOI221_X1 port map( B1 => n2562, B2 => n3142, C1 => n2563, C2 => 
                           n3133, A => n2692, ZN => n2689);
   U2440 : OAI22_X1 port map( A1 => n1821, A2 => n2565, B1 => n1861, B2 => 
                           n2566, ZN => n2692);
   U2441 : AOI21_X1 port map( B1 => n2693, B2 => n2694, A => n2574, ZN => n2682
                           );
   U2442 : OAI22_X1 port map( A1 => n1899, A2 => n2560, B1 => n3131, B2 => 
                           n2561, ZN => n2695);
   U2443 : OAI22_X1 port map( A1 => n1962, A2 => n2565, B1 => n1869, B2 => 
                           n2566, ZN => n2696);
   U2444 : AOI21_X1 port map( B1 => n2697, B2 => n2698, A => n2579, ZN => n2681
                           );
   U2445 : OAI22_X1 port map( A1 => n3134, A2 => n2560, B1 => n1836, B2 => 
                           n2561, ZN => n2699);
   U2446 : OAI22_X1 port map( A1 => n1963, A2 => n2565, B1 => n1805, B2 => 
                           n2566, ZN => n2700);
   U2447 : OAI22_X1 port map( A1 => n3042, A2 => n2585, B1 => n1923, B2 => 
                           n2586, ZN => n2701);
   U2448 : NAND2_X1 port map( A1 => n2702, A2 => n2703, ZN => n1258);
   U2449 : NOR4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => n2707
                           , ZN => n2703);
   U2450 : AOI21_X1 port map( B1 => n2708, B2 => n2709, A => n2556, ZN => n2707
                           );
   U2451 : INV_X1 port map( A => n2710, ZN => n2556);
   U2452 : OAI22_X1 port map( A1 => n3123, A2 => n2560, B1 => n1814, B2 => 
                           n2561, ZN => n2711);
   U2453 : OAI22_X1 port map( A1 => n1972, A2 => n2565, B1 => n1862, B2 => 
                           n2566, ZN => n2712);
   U2454 : AOI21_X1 port map( B1 => n2713, B2 => n2714, A => n2569, ZN => n2706
                           );
   U2455 : INV_X1 port map( A => n2715, ZN => n2569);
   U2456 : OAI22_X1 port map( A1 => n3124, A2 => n2560, B1 => n3035, B2 => 
                           n2561, ZN => n2716);
   U2457 : OAI22_X1 port map( A1 => n1822, A2 => n2565, B1 => n1863, B2 => 
                           n2566, ZN => n2717);
   U2458 : AOI21_X1 port map( B1 => n2718, B2 => n2719, A => n2574, ZN => n2705
                           );
   U2459 : OAI22_X1 port map( A1 => n1900, A2 => n2560, B1 => n3119, B2 => 
                           n2561, ZN => n2720);
   U2460 : OAI22_X1 port map( A1 => n1964, A2 => n2565, B1 => n1870, B2 => 
                           n2566, ZN => n2721);
   U2461 : AOI21_X1 port map( B1 => n2722, B2 => n2723, A => n2579, ZN => n2704
                           );
   U2462 : OAI22_X1 port map( A1 => n3122, A2 => n2560, B1 => n1837, B2 => 
                           n2561, ZN => n2724);
   U2463 : OAI22_X1 port map( A1 => n1965, A2 => n2565, B1 => n1806, B2 => 
                           n2566, ZN => n2725);
   U2464 : OAI22_X1 port map( A1 => n3043, A2 => n2585, B1 => n1924, B2 => 
                           n2586, ZN => n2726);
   U2465 : NAND2_X1 port map( A1 => RD2, A2 => n2727, ZN => n1257);
   U2466 : NAND4_X1 port map( A1 => n2728, A2 => n2729, A3 => n2730, A4 => 
                           n2731, ZN => n1256);
   U2467 : INV_X1 port map( A => n2732, ZN => n2731);
   U2468 : OAI221_X1 port map( B1 => n2586, B2 => n1933, C1 => n2585, C2 => 
                           n3044, A => n2733, ZN => n2732);
   U2469 : INV_X1 port map( A => n2734, ZN => n2733);
   U2470 : OAI22_X1 port map( A1 => n2735, A2 => n2574, B1 => n2736, B2 => 
                           n2579, ZN => n2734);
   U2471 : NAND3_X1 port map( A1 => n2737, A2 => n2738, A3 => n2739, ZN => 
                           n2579);
   U2472 : NOR4_X1 port map( A1 => n2740, A2 => n2741, A3 => n2742, A4 => n2743
                           , ZN => n2736);
   U2473 : OAI22_X1 port map( A1 => n1848, A2 => n2565, B1 => n1890, B2 => 
                           n2566, ZN => n2743);
   U2474 : OAI22_X1 port map( A1 => n1815, A2 => n2744, B1 => n1908, B2 => 
                           n2745, ZN => n2742);
   U2475 : OAI22_X1 port map( A1 => n3112, A2 => n2560, B1 => n1838, B2 => 
                           n2561, ZN => n2741);
   U2476 : OAI22_X1 port map( A1 => n1807, A2 => n2746, B1 => n3222, B2 => 
                           n2747, ZN => n2740);
   U2477 : NAND3_X1 port map( A1 => n2748, A2 => n2738, A3 => n2737, ZN => 
                           n2574);
   U2478 : NOR4_X1 port map( A1 => n2749, A2 => n2750, A3 => n2751, A4 => n2752
                           , ZN => n2735);
   U2479 : OAI22_X1 port map( A1 => n1849, A2 => n2565, B1 => n1910, B2 => 
                           n2566, ZN => n2752);
   U2480 : OAI22_X1 port map( A1 => n1839, A2 => n2744, B1 => n1909, B2 => 
                           n2745, ZN => n2751);
   U2481 : OAI22_X1 port map( A1 => n1901, A2 => n2560, B1 => n3109, B2 => 
                           n2561, ZN => n2750);
   U2482 : OAI22_X1 port map( A1 => n1907, A2 => n2746, B1 => n1799, B2 => 
                           n2747, ZN => n2749);
   U2483 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => n2753, A3 => n2754, ZN =>
                           n2585);
   U2484 : NAND3_X1 port map( A1 => n2753, A2 => n2755, A3 => n2754, ZN => 
                           n2586);
   U2485 : AOI22_X1 port map( A1 => n2582, A2 => n1936, B1 => n2583, B2 => 
                           n3101, ZN => n2730);
   U2486 : OAI21_X1 port map( B1 => n2756, B2 => n2757, A => n2715, ZN => n2729
                           );
   U2487 : NOR3_X1 port map( A1 => n2739, A2 => n2754, A3 => n2737, ZN => n2715
                           );
   U2488 : OAI221_X1 port map( B1 => n1932, B2 => n2566, C1 => n1880, C2 => 
                           n2565, A => n2758, ZN => n2757);
   U2489 : AOI22_X1 port map( A1 => n2562, A2 => n3118, B1 => n2563, B2 => 
                           n3111, ZN => n2758);
   U2490 : OAI221_X1 port map( B1 => n3036, B2 => n2561, C1 => n3114, C2 => 
                           n2560, A => n2759, ZN => n2756);
   U2491 : AOI22_X1 port map( A1 => n2557, A2 => n1935, B1 => n2558, B2 => 
                           n3115, ZN => n2759);
   U2492 : OAI21_X1 port map( B1 => n2760, B2 => n2761, A => n2710, ZN => n2728
                           );
   U2493 : NOR3_X1 port map( A1 => n2737, A2 => n2754, A3 => n2748, ZN => n2710
                           );
   U2494 : INV_X1 port map( A => n2739, ZN => n2748);
   U2495 : XNOR2_X1 port map( A => n2762, B => n2763, ZN => n2739);
   U2496 : XOR2_X1 port map( A => ADD_RD2(2), B => CWP_2_port, Z => n2762);
   U2497 : INV_X1 port map( A => n2738, ZN => n2754);
   U2498 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(2), ZN => n2738);
   U2499 : XNOR2_X1 port map( A => n2764, B => n2765, ZN => n2737);
   U2500 : XOR2_X1 port map( A => n1489, B => ADD_RD2(1), Z => n2765);
   U2501 : OAI221_X1 port map( B1 => n1872, B2 => n2566, C1 => n1996, C2 => 
                           n2565, A => n2766, ZN => n2761);
   U2502 : AOI22_X1 port map( A1 => n2562, A2 => n3053, B1 => n2563, B2 => 
                           n3110, ZN => n2766);
   U2503 : NAND3_X1 port map( A1 => n2767, A2 => n2768, A3 => n2769, ZN => 
                           n2744);
   U2504 : NAND3_X1 port map( A1 => n2770, A2 => n2768, A3 => n2767, ZN => 
                           n2745);
   U2505 : INV_X1 port map( A => n2772, ZN => n2768);
   U2506 : OAI221_X1 port map( B1 => n1891, B2 => n2561, C1 => n3113, C2 => 
                           n2560, A => n2773, ZN => n2760);
   U2507 : AOI22_X1 port map( A1 => n2557, A2 => n1840, B1 => n2558, B2 => 
                           n3116, ZN => n2773);
   U2508 : NAND3_X1 port map( A1 => n2772, A2 => n2770, A3 => n2767, ZN => 
                           n2746);
   U2509 : NAND3_X1 port map( A1 => n2770, A2 => n2771, A3 => n2772, ZN => 
                           n2747);
   U2510 : INV_X1 port map( A => n2770, ZN => n2769);
   U2511 : XOR2_X1 port map( A => n1490, B => ADD_RD2(0), Z => n2770);
   U2512 : INV_X1 port map( A => n2767, ZN => n2771);
   U2513 : XNOR2_X1 port map( A => n2774, B => n2775, ZN => n2767);
   U2514 : XOR2_X1 port map( A => n1487, B => ADD_RD2(3), Z => n2775);
   U2515 : XOR2_X1 port map( A => n2776, B => n1486, Z => n2772);
   U2516 : OAI22_X1 port map( A1 => n2774, A2 => n2777, B1 => n1487, B2 => 
                           n2778, ZN => n2776);
   U2517 : AND2_X1 port map( A1 => n2777, A2 => n2774, ZN => n2778);
   U2518 : INV_X1 port map( A => ADD_RD2(3), ZN => n2777);
   U2519 : AOI21_X1 port map( B1 => n2763, B2 => ADD_RD2(2), A => n2779, ZN => 
                           n2774);
   U2520 : INV_X1 port map( A => n2780, ZN => n2779);
   U2521 : OAI21_X1 port map( B1 => ADD_RD2(2), B2 => n2763, A => CWP_2_port, 
                           ZN => n2780);
   U2522 : OAI21_X1 port map( B1 => n2781, B2 => n2755, A => n2782, ZN => n2763
                           );
   U2523 : INV_X1 port map( A => n2783, ZN => n2782);
   U2524 : AOI21_X1 port map( B1 => n2781, B2 => n2755, A => n1489, ZN => n2783
                           );
   U2525 : INV_X1 port map( A => ADD_RD2(1), ZN => n2755);
   U2526 : INV_X1 port map( A => n2764, ZN => n2781);
   U2527 : NOR2_X1 port map( A1 => n2753, A2 => n1490, ZN => n2764);
   U2528 : INV_X1 port map( A => ADD_RD2(0), ZN => n2753);
   U2529 : NAND2_X1 port map( A1 => n2784, A2 => n2785, ZN => n1255);
   U2530 : NOR4_X1 port map( A1 => n2786, A2 => n2787, A3 => n2788, A4 => n2789
                           , ZN => n2785);
   U2531 : AOI21_X1 port map( B1 => n2790, B2 => n2791, A => n2792, ZN => n2789
                           );
   U2532 : AOI221_X1 port map( B1 => n2043, B2 => n1842, C1 => n2045, C2 => 
                           n3198, A => n2795, ZN => n2791);
   U2533 : OAI22_X1 port map( A1 => n3195, A2 => n2796, B1 => n1808, B2 => 
                           n2797, ZN => n2795);
   U2534 : AOI221_X1 port map( B1 => n2044, B2 => n3060, C1 => n2046, C2 => 
                           n3084, A => n2800, ZN => n2790);
   U2535 : OAI22_X1 port map( A1 => n1850, A2 => n2801, B1 => n1973, B2 => 
                           n2802, ZN => n2800);
   U2536 : AOI21_X1 port map( B1 => n2803, B2 => n2804, A => n2805, ZN => n2788
                           );
   U2537 : AOI221_X1 port map( B1 => n2043, B2 => n1938, C1 => n2045, C2 => 
                           n3197, A => n2806, ZN => n2804);
   U2538 : OAI22_X1 port map( A1 => n3196, A2 => n2796, B1 => n3029, B2 => 
                           n2797, ZN => n2806);
   U2539 : AOI221_X1 port map( B1 => n2044, B2 => n3202, C1 => n2046, C2 => 
                           n3201, A => n2807, ZN => n2803);
   U2540 : OAI22_X1 port map( A1 => n1851, A2 => n2801, B1 => n1911, B2 => 
                           n2802, ZN => n2807);
   U2541 : AOI21_X1 port map( B1 => n2808, B2 => n2809, A => n2810, ZN => n2787
                           );
   U2542 : AOI221_X1 port map( B1 => n2043, B2 => n3200, C1 => n2045, C2 => 
                           n3052, A => n2811, ZN => n2809);
   U2543 : OAI22_X1 port map( A1 => n1894, A2 => n2796, B1 => n3191, B2 => 
                           n2797, ZN => n2811);
   U2544 : AOI221_X1 port map( B1 => n2044, B2 => n3076, C1 => n2046, C2 => 
                           n3218, A => n2812, ZN => n2808);
   U2545 : OAI22_X1 port map( A1 => n1864, A2 => n2801, B1 => n1925, B2 => 
                           n2802, ZN => n2812);
   U2546 : AOI21_X1 port map( B1 => n2813, B2 => n2814, A => n2815, ZN => n2786
                           );
   U2547 : AOI221_X1 port map( B1 => n2043, B2 => n1902, C1 => n2045, C2 => 
                           n3199, A => n2816, ZN => n2814);
   U2548 : OAI22_X1 port map( A1 => n3194, A2 => n2796, B1 => n1831, B2 => 
                           n2797, ZN => n2816);
   U2549 : AOI221_X1 port map( B1 => n2044, B2 => n3068, C1 => n2046, C2 => 
                           n3217, A => n2817, ZN => n2813);
   U2550 : OAI22_X1 port map( A1 => n1800, A2 => n2801, B1 => n1873, B2 => 
                           n2802, ZN => n2817);
   U2551 : AOI221_X1 port map( B1 => n2818, B2 => n1951, C1 => n2819, C2 => 
                           n3108, A => n2820, ZN => n2784);
   U2552 : OAI22_X1 port map( A1 => n3037, A2 => n2821, B1 => n1918, B2 => 
                           n2822, ZN => n2820);
   U2553 : NAND2_X1 port map( A1 => n2823, A2 => n2824, ZN => n1254);
   U2554 : NOR4_X1 port map( A1 => n2825, A2 => n2826, A3 => n2827, A4 => n2828
                           , ZN => n2824);
   U2555 : AOI21_X1 port map( B1 => n2829, B2 => n2830, A => n2792, ZN => n2828
                           );
   U2556 : AOI221_X1 port map( B1 => n2043, B2 => n1843, C1 => n2045, C2 => 
                           n3186, A => n2831, ZN => n2830);
   U2557 : OAI22_X1 port map( A1 => n3183, A2 => n2796, B1 => n1809, B2 => 
                           n2797, ZN => n2831);
   U2558 : AOI221_X1 port map( B1 => n2044, B2 => n3059, C1 => n2046, C2 => 
                           n3083, A => n2832, ZN => n2829);
   U2559 : OAI22_X1 port map( A1 => n1852, A2 => n2801, B1 => n1974, B2 => 
                           n2802, ZN => n2832);
   U2560 : AOI21_X1 port map( B1 => n2833, B2 => n2834, A => n2805, ZN => n2827
                           );
   U2561 : AOI221_X1 port map( B1 => n2043, B2 => n1939, C1 => n2045, C2 => 
                           n3185, A => n2835, ZN => n2834);
   U2562 : OAI22_X1 port map( A1 => n3184, A2 => n2796, B1 => n3030, B2 => 
                           n2797, ZN => n2835);
   U2563 : AOI221_X1 port map( B1 => n2044, B2 => n3190, C1 => n2046, C2 => 
                           n3189, A => n2836, ZN => n2833);
   U2564 : OAI22_X1 port map( A1 => n1853, A2 => n2801, B1 => n1912, B2 => 
                           n2802, ZN => n2836);
   U2565 : AOI21_X1 port map( B1 => n2837, B2 => n2838, A => n2810, ZN => n2826
                           );
   U2566 : AOI221_X1 port map( B1 => n2043, B2 => n3188, C1 => n2045, C2 => 
                           n3051, A => n2839, ZN => n2838);
   U2567 : OAI22_X1 port map( A1 => n1895, A2 => n2796, B1 => n3179, B2 => 
                           n2797, ZN => n2839);
   U2568 : AOI221_X1 port map( B1 => n2044, B2 => n3075, C1 => n2046, C2 => 
                           n3216, A => n2840, ZN => n2837);
   U2569 : OAI22_X1 port map( A1 => n1865, A2 => n2801, B1 => n1926, B2 => 
                           n2802, ZN => n2840);
   U2570 : AOI21_X1 port map( B1 => n2841, B2 => n2842, A => n2815, ZN => n2825
                           );
   U2571 : AOI221_X1 port map( B1 => n2043, B2 => n1903, C1 => n2045, C2 => 
                           n3187, A => n2843, ZN => n2842);
   U2572 : OAI22_X1 port map( A1 => n3182, A2 => n2796, B1 => n1832, B2 => 
                           n2797, ZN => n2843);
   U2573 : AOI221_X1 port map( B1 => n2044, B2 => n3067, C1 => n2046, C2 => 
                           n3215, A => n2844, ZN => n2841);
   U2574 : OAI22_X1 port map( A1 => n1801, A2 => n2801, B1 => n1874, B2 => 
                           n2802, ZN => n2844);
   U2575 : OAI22_X1 port map( A1 => n3038, A2 => n2821, B1 => n1919, B2 => 
                           n2822, ZN => n2845);
   U2576 : NAND2_X1 port map( A1 => n2846, A2 => n2847, ZN => n1253);
   U2577 : NOR4_X1 port map( A1 => n2848, A2 => n2849, A3 => n2850, A4 => n2851
                           , ZN => n2847);
   U2578 : AOI21_X1 port map( B1 => n2852, B2 => n2853, A => n2792, ZN => n2851
                           );
   U2579 : AOI221_X1 port map( B1 => n2043, B2 => n1844, C1 => n2045, C2 => 
                           n3174, A => n2854, ZN => n2853);
   U2580 : OAI22_X1 port map( A1 => n3171, A2 => n2796, B1 => n1810, B2 => 
                           n2797, ZN => n2854);
   U2581 : AOI221_X1 port map( B1 => n2044, B2 => n3058, C1 => n2046, C2 => 
                           n3082, A => n2855, ZN => n2852);
   U2582 : OAI22_X1 port map( A1 => n1854, A2 => n2801, B1 => n1975, B2 => 
                           n2802, ZN => n2855);
   U2583 : AOI21_X1 port map( B1 => n2856, B2 => n2857, A => n2805, ZN => n2850
                           );
   U2584 : AOI221_X1 port map( B1 => n2043, B2 => n1940, C1 => n2045, C2 => 
                           n3173, A => n2858, ZN => n2857);
   U2585 : OAI22_X1 port map( A1 => n3172, A2 => n2796, B1 => n3031, B2 => 
                           n2797, ZN => n2858);
   U2586 : AOI221_X1 port map( B1 => n2044, B2 => n3178, C1 => n2046, C2 => 
                           n3177, A => n2859, ZN => n2856);
   U2587 : OAI22_X1 port map( A1 => n1855, A2 => n2801, B1 => n1913, B2 => 
                           n2802, ZN => n2859);
   U2588 : AOI21_X1 port map( B1 => n2860, B2 => n2861, A => n2810, ZN => n2849
                           );
   U2589 : AOI221_X1 port map( B1 => n2043, B2 => n3176, C1 => n2045, C2 => 
                           n3050, A => n2862, ZN => n2861);
   U2590 : OAI22_X1 port map( A1 => n1896, A2 => n2796, B1 => n3167, B2 => 
                           n2797, ZN => n2862);
   U2591 : AOI221_X1 port map( B1 => n2044, B2 => n3074, C1 => n2046, C2 => 
                           n3214, A => n2863, ZN => n2860);
   U2592 : OAI22_X1 port map( A1 => n1866, A2 => n2801, B1 => n1927, B2 => 
                           n2802, ZN => n2863);
   U2593 : AOI21_X1 port map( B1 => n2864, B2 => n2865, A => n2815, ZN => n2848
                           );
   U2594 : AOI221_X1 port map( B1 => n2043, B2 => n1904, C1 => n2045, C2 => 
                           n3175, A => n2866, ZN => n2865);
   U2595 : OAI22_X1 port map( A1 => n3170, A2 => n2796, B1 => n1833, B2 => 
                           n2797, ZN => n2866);
   U2596 : AOI221_X1 port map( B1 => n2044, B2 => n3066, C1 => n2046, C2 => 
                           n3213, A => n2867, ZN => n2864);
   U2597 : OAI22_X1 port map( A1 => n1802, A2 => n2801, B1 => n1875, B2 => 
                           n2802, ZN => n2867);
   U2598 : OAI22_X1 port map( A1 => n3039, A2 => n2821, B1 => n1920, B2 => 
                           n2822, ZN => n2868);
   U2599 : NAND2_X1 port map( A1 => n2869, A2 => n2870, ZN => n1252);
   U2600 : NOR4_X1 port map( A1 => n2871, A2 => n2872, A3 => n2873, A4 => n2874
                           , ZN => n2870);
   U2601 : AOI21_X1 port map( B1 => n2875, B2 => n2876, A => n2792, ZN => n2874
                           );
   U2602 : AOI221_X1 port map( B1 => n2043, B2 => n1845, C1 => n2045, C2 => 
                           n3162, A => n2877, ZN => n2876);
   U2603 : OAI22_X1 port map( A1 => n3159, A2 => n2796, B1 => n1811, B2 => 
                           n2797, ZN => n2877);
   U2604 : AOI221_X1 port map( B1 => n2044, B2 => n3057, C1 => n2046, C2 => 
                           n3081, A => n2878, ZN => n2875);
   U2605 : OAI22_X1 port map( A1 => n1856, A2 => n2801, B1 => n1976, B2 => 
                           n2802, ZN => n2878);
   U2606 : AOI21_X1 port map( B1 => n2879, B2 => n2880, A => n2805, ZN => n2873
                           );
   U2607 : AOI221_X1 port map( B1 => n2043, B2 => n1941, C1 => n2045, C2 => 
                           n3161, A => n2881, ZN => n2880);
   U2608 : OAI22_X1 port map( A1 => n3160, A2 => n2796, B1 => n3032, B2 => 
                           n2797, ZN => n2881);
   U2609 : AOI221_X1 port map( B1 => n2044, B2 => n3166, C1 => n2046, C2 => 
                           n3165, A => n2882, ZN => n2879);
   U2610 : OAI22_X1 port map( A1 => n1857, A2 => n2801, B1 => n1914, B2 => 
                           n2802, ZN => n2882);
   U2611 : AOI21_X1 port map( B1 => n2883, B2 => n2884, A => n2810, ZN => n2872
                           );
   U2612 : AOI221_X1 port map( B1 => n2043, B2 => n3164, C1 => n2045, C2 => 
                           n3049, A => n2885, ZN => n2884);
   U2613 : OAI22_X1 port map( A1 => n1897, A2 => n2796, B1 => n3155, B2 => 
                           n2797, ZN => n2885);
   U2614 : AOI221_X1 port map( B1 => n2044, B2 => n3073, C1 => n2046, C2 => 
                           n3212, A => n2886, ZN => n2883);
   U2615 : OAI22_X1 port map( A1 => n1867, A2 => n2801, B1 => n1928, B2 => 
                           n2802, ZN => n2886);
   U2616 : AOI21_X1 port map( B1 => n2887, B2 => n2888, A => n2815, ZN => n2871
                           );
   U2617 : AOI221_X1 port map( B1 => n2043, B2 => n1905, C1 => n2045, C2 => 
                           n3163, A => n2889, ZN => n2888);
   U2618 : OAI22_X1 port map( A1 => n3158, A2 => n2796, B1 => n1834, B2 => 
                           n2797, ZN => n2889);
   U2619 : AOI221_X1 port map( B1 => n2044, B2 => n3065, C1 => n2046, C2 => 
                           n3211, A => n2890, ZN => n2887);
   U2620 : OAI22_X1 port map( A1 => n1803, A2 => n2801, B1 => n1876, B2 => 
                           n2802, ZN => n2890);
   U2621 : OAI22_X1 port map( A1 => n3040, A2 => n2821, B1 => n1921, B2 => 
                           n2822, ZN => n2891);
   U2622 : NAND2_X1 port map( A1 => n2892, A2 => n2893, ZN => n1251);
   U2623 : NOR4_X1 port map( A1 => n2894, A2 => n2895, A3 => n2896, A4 => n2897
                           , ZN => n2893);
   U2624 : AOI21_X1 port map( B1 => n2898, B2 => n2899, A => n2792, ZN => n2897
                           );
   U2625 : AOI221_X1 port map( B1 => n2043, B2 => n1846, C1 => n2045, C2 => 
                           n3150, A => n2900, ZN => n2899);
   U2626 : OAI22_X1 port map( A1 => n3147, A2 => n2796, B1 => n1812, B2 => 
                           n2797, ZN => n2900);
   U2627 : AOI221_X1 port map( B1 => n2044, B2 => n3056, C1 => n2046, C2 => 
                           n3080, A => n2901, ZN => n2898);
   U2628 : OAI22_X1 port map( A1 => n1858, A2 => n2801, B1 => n1977, B2 => 
                           n2802, ZN => n2901);
   U2629 : AOI21_X1 port map( B1 => n2902, B2 => n2903, A => n2805, ZN => n2896
                           );
   U2630 : AOI221_X1 port map( B1 => n2043, B2 => n1942, C1 => n2045, C2 => 
                           n3149, A => n2904, ZN => n2903);
   U2631 : OAI22_X1 port map( A1 => n3148, A2 => n2796, B1 => n3033, B2 => 
                           n2797, ZN => n2904);
   U2632 : AOI221_X1 port map( B1 => n2044, B2 => n3154, C1 => n2046, C2 => 
                           n3153, A => n2905, ZN => n2902);
   U2633 : OAI22_X1 port map( A1 => n1859, A2 => n2801, B1 => n1915, B2 => 
                           n2802, ZN => n2905);
   U2634 : AOI21_X1 port map( B1 => n2906, B2 => n2907, A => n2810, ZN => n2895
                           );
   U2635 : AOI221_X1 port map( B1 => n2043, B2 => n3152, C1 => n2045, C2 => 
                           n3048, A => n2908, ZN => n2907);
   U2636 : OAI22_X1 port map( A1 => n1898, A2 => n2796, B1 => n3143, B2 => 
                           n2797, ZN => n2908);
   U2637 : AOI221_X1 port map( B1 => n2044, B2 => n3072, C1 => n2046, C2 => 
                           n3210, A => n2909, ZN => n2906);
   U2638 : OAI22_X1 port map( A1 => n1868, A2 => n2801, B1 => n1929, B2 => 
                           n2802, ZN => n2909);
   U2639 : AOI21_X1 port map( B1 => n2910, B2 => n2911, A => n2815, ZN => n2894
                           );
   U2640 : AOI221_X1 port map( B1 => n2043, B2 => n1906, C1 => n2045, C2 => 
                           n3151, A => n2912, ZN => n2911);
   U2641 : OAI22_X1 port map( A1 => n3146, A2 => n2796, B1 => n1835, B2 => 
                           n2797, ZN => n2912);
   U2642 : AOI221_X1 port map( B1 => n2044, B2 => n3064, C1 => n2046, C2 => 
                           n3209, A => n2913, ZN => n2910);
   U2643 : OAI22_X1 port map( A1 => n1804, A2 => n2801, B1 => n1877, B2 => 
                           n2802, ZN => n2913);
   U2644 : OAI22_X1 port map( A1 => n3041, A2 => n2821, B1 => n1922, B2 => 
                           n2822, ZN => n2914);
   U2645 : NAND2_X1 port map( A1 => n2915, A2 => n2916, ZN => n1250);
   U2646 : NOR4_X1 port map( A1 => n2917, A2 => n2918, A3 => n2919, A4 => n2920
                           , ZN => n2916);
   U2647 : AOI21_X1 port map( B1 => n2921, B2 => n2922, A => n2792, ZN => n2920
                           );
   U2648 : AOI221_X1 port map( B1 => n2043, B2 => n1847, C1 => n2045, C2 => 
                           n3138, A => n2923, ZN => n2922);
   U2649 : OAI22_X1 port map( A1 => n3135, A2 => n2796, B1 => n1813, B2 => 
                           n2797, ZN => n2923);
   U2650 : AOI221_X1 port map( B1 => n2044, B2 => n3055, C1 => n2046, C2 => 
                           n3079, A => n2924, ZN => n2921);
   U2651 : OAI22_X1 port map( A1 => n1860, A2 => n2801, B1 => n1978, B2 => 
                           n2802, ZN => n2924);
   U2652 : AOI21_X1 port map( B1 => n2925, B2 => n2926, A => n2805, ZN => n2919
                           );
   U2653 : AOI221_X1 port map( B1 => n2043, B2 => n1943, C1 => n2045, C2 => 
                           n3137, A => n2927, ZN => n2926);
   U2654 : OAI22_X1 port map( A1 => n3136, A2 => n2796, B1 => n3034, B2 => 
                           n2797, ZN => n2927);
   U2655 : AOI221_X1 port map( B1 => n2044, B2 => n3142, C1 => n2046, C2 => 
                           n3141, A => n2928, ZN => n2925);
   U2656 : OAI22_X1 port map( A1 => n1861, A2 => n2801, B1 => n1916, B2 => 
                           n2802, ZN => n2928);
   U2657 : AOI21_X1 port map( B1 => n2929, B2 => n2930, A => n2810, ZN => n2918
                           );
   U2658 : AOI221_X1 port map( B1 => n2043, B2 => n3140, C1 => n2794, C2 => 
                           n3047, A => n2931, ZN => n2930);
   U2659 : OAI22_X1 port map( A1 => n1899, A2 => n2796, B1 => n3131, B2 => 
                           n2797, ZN => n2931);
   U2660 : AOI221_X1 port map( B1 => n2044, B2 => n3071, C1 => n2799, C2 => 
                           n3208, A => n2932, ZN => n2929);
   U2661 : OAI22_X1 port map( A1 => n1869, A2 => n2801, B1 => n1930, B2 => 
                           n2802, ZN => n2932);
   U2662 : AOI21_X1 port map( B1 => n2933, B2 => n2934, A => n2815, ZN => n2917
                           );
   U2663 : AOI221_X1 port map( B1 => n2043, B2 => n1892, C1 => n2794, C2 => 
                           n3139, A => n2935, ZN => n2934);
   U2664 : OAI22_X1 port map( A1 => n3134, A2 => n2796, B1 => n1836, B2 => 
                           n2797, ZN => n2935);
   U2665 : AOI221_X1 port map( B1 => n2044, B2 => n3063, C1 => n2799, C2 => 
                           n3207, A => n2936, ZN => n2933);
   U2666 : OAI22_X1 port map( A1 => n1805, A2 => n2801, B1 => n1878, B2 => 
                           n2802, ZN => n2936);
   U2667 : OAI22_X1 port map( A1 => n3042, A2 => n2821, B1 => n1923, B2 => 
                           n2822, ZN => n2937);
   U2668 : NAND2_X1 port map( A1 => n2938, A2 => n2939, ZN => n1249);
   U2669 : NOR4_X1 port map( A1 => n2940, A2 => n2941, A3 => n2942, A4 => n2943
                           , ZN => n2939);
   U2670 : AOI21_X1 port map( B1 => n2944, B2 => n2945, A => n2792, ZN => n2943
                           );
   U2671 : INV_X1 port map( A => n2946, ZN => n2792);
   U2672 : AOI221_X1 port map( B1 => n2793, B2 => n1841, C1 => n2794, C2 => 
                           n3126, A => n2947, ZN => n2945);
   U2673 : OAI22_X1 port map( A1 => n3123, A2 => n2796, B1 => n1814, B2 => 
                           n2797, ZN => n2947);
   U2674 : AOI221_X1 port map( B1 => n2798, B2 => n3054, C1 => n2799, C2 => 
                           n3078, A => n2948, ZN => n2944);
   U2675 : OAI22_X1 port map( A1 => n1862, A2 => n2801, B1 => n1979, B2 => 
                           n2802, ZN => n2948);
   U2676 : AOI21_X1 port map( B1 => n2949, B2 => n2950, A => n2805, ZN => n2942
                           );
   U2677 : INV_X1 port map( A => n2951, ZN => n2805);
   U2678 : AOI221_X1 port map( B1 => n2793, B2 => n1937, C1 => n2794, C2 => 
                           n3125, A => n2952, ZN => n2950);
   U2679 : OAI22_X1 port map( A1 => n3124, A2 => n2796, B1 => n3035, B2 => 
                           n2797, ZN => n2952);
   U2680 : AOI221_X1 port map( B1 => n2798, B2 => n3130, C1 => n2799, C2 => 
                           n3129, A => n2953, ZN => n2949);
   U2681 : OAI22_X1 port map( A1 => n1863, A2 => n2801, B1 => n1917, B2 => 
                           n2802, ZN => n2953);
   U2682 : AOI21_X1 port map( B1 => n2954, B2 => n2955, A => n2810, ZN => n2941
                           );
   U2683 : AOI221_X1 port map( B1 => n2793, B2 => n3128, C1 => n2794, C2 => 
                           n3046, A => n2956, ZN => n2955);
   U2684 : OAI22_X1 port map( A1 => n1900, A2 => n2796, B1 => n3119, B2 => 
                           n2797, ZN => n2956);
   U2685 : AOI221_X1 port map( B1 => n2798, B2 => n3070, C1 => n2799, C2 => 
                           n3206, A => n2957, ZN => n2954);
   U2686 : OAI22_X1 port map( A1 => n1870, A2 => n2801, B1 => n1931, B2 => 
                           n2802, ZN => n2957);
   U2687 : AOI21_X1 port map( B1 => n2958, B2 => n2959, A => n2815, ZN => n2940
                           );
   U2688 : AOI221_X1 port map( B1 => n2793, B2 => n1893, C1 => n2794, C2 => 
                           n3127, A => n2960, ZN => n2959);
   U2689 : OAI22_X1 port map( A1 => n3122, A2 => n2796, B1 => n1837, B2 => 
                           n2797, ZN => n2960);
   U2690 : AOI221_X1 port map( B1 => n2798, B2 => n3062, C1 => n2799, C2 => 
                           n3205, A => n2961, ZN => n2958);
   U2691 : OAI22_X1 port map( A1 => n1806, A2 => n2801, B1 => n1879, B2 => 
                           n2802, ZN => n2961);
   U2692 : OAI22_X1 port map( A1 => n3043, A2 => n2821, B1 => n1924, B2 => 
                           n2822, ZN => n2962);
   U2693 : NAND2_X1 port map( A1 => RD1, A2 => n2727, ZN => n1248);
   U2694 : AND4_X1 port map( A1 => ENABLE, A2 => n2139, A3 => n2144, A4 => 
                           n2142, ZN => n2727);
   U2695 : NOR2_X1 port map( A1 => n3286, A2 => SPILL_port, ZN => n2139);
   U2696 : INV_X1 port map( A => n1266, ZN => SPILL_port);
   U2697 : NAND4_X1 port map( A1 => n2963, A2 => n2964, A3 => n2965, A4 => 
                           n2966, ZN => n1247);
   U2698 : INV_X1 port map( A => n2967, ZN => n2966);
   U2699 : OAI221_X1 port map( B1 => n2822, B2 => n1933, C1 => n2821, C2 => 
                           n3044, A => n2968, ZN => n2967);
   U2700 : INV_X1 port map( A => n2969, ZN => n2968);
   U2701 : OAI22_X1 port map( A1 => n2970, A2 => n2810, B1 => n2971, B2 => 
                           n2815, ZN => n2969);
   U2702 : NAND3_X1 port map( A1 => n2972, A2 => n2973, A3 => n2974, ZN => 
                           n2815);
   U2703 : NOR4_X1 port map( A1 => n2975, A2 => n2976, A3 => n2977, A4 => n2978
                           , ZN => n2971);
   U2704 : OAI22_X1 port map( A1 => n1890, A2 => n2801, B1 => n1815, B2 => 
                           n2802, ZN => n2978);
   U2705 : OAI22_X1 port map( A1 => n1848, A2 => n2979, B1 => n1908, B2 => 
                           n2980, ZN => n2977);
   U2706 : OAI22_X1 port map( A1 => n3112, A2 => n2796, B1 => n1838, B2 => 
                           n2797, ZN => n2976);
   U2707 : OAI22_X1 port map( A1 => n1807, A2 => n2981, B1 => n3222, B2 => 
                           n2982, ZN => n2975);
   U2708 : NAND3_X1 port map( A1 => n2983, A2 => n2973, A3 => n2972, ZN => 
                           n2810);
   U2709 : NOR4_X1 port map( A1 => n2984, A2 => n2985, A3 => n2986, A4 => n2987
                           , ZN => n2970);
   U2710 : OAI22_X1 port map( A1 => n1910, A2 => n2801, B1 => n1839, B2 => 
                           n2802, ZN => n2987);
   U2711 : OAI22_X1 port map( A1 => n1849, A2 => n2979, B1 => n1909, B2 => 
                           n2980, ZN => n2986);
   U2712 : INV_X1 port map( A => n2798, ZN => n2980);
   U2713 : INV_X1 port map( A => n2799, ZN => n2979);
   U2714 : OAI22_X1 port map( A1 => n1901, A2 => n2796, B1 => n3109, B2 => 
                           n2797, ZN => n2985);
   U2715 : OAI22_X1 port map( A1 => n1907, A2 => n2981, B1 => n1799, B2 => 
                           n2982, ZN => n2984);
   U2716 : INV_X1 port map( A => n2793, ZN => n2982);
   U2717 : INV_X1 port map( A => n2794, ZN => n2981);
   U2718 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => n2988, A3 => n2989, ZN =>
                           n2821);
   U2719 : NAND3_X1 port map( A1 => n2988, A2 => n2990, A3 => n2989, ZN => 
                           n2822);
   U2720 : AOI22_X1 port map( A1 => n2818, A2 => n1936, B1 => n2819, B2 => 
                           n3101, ZN => n2965);
   U2721 : OAI21_X1 port map( B1 => n2991, B2 => n2992, A => n2951, ZN => n2964
                           );
   U2722 : NOR3_X1 port map( A1 => n2974, A2 => n2989, A3 => n2972, ZN => n2951
                           );
   U2723 : OAI221_X1 port map( B1 => n1871, B2 => n2802, C1 => n1932, C2 => 
                           n2801, A => n2993, ZN => n2992);
   U2724 : AOI22_X1 port map( A1 => n2798, A2 => n3118, B1 => n2046, B2 => 
                           n3117, ZN => n2993);
   U2725 : OAI221_X1 port map( B1 => n3036, B2 => n2797, C1 => n3114, C2 => 
                           n2796, A => n2994, ZN => n2991);
   U2726 : AOI22_X1 port map( A1 => n2793, A2 => n1935, B1 => n2045, B2 => 
                           n3115, ZN => n2994);
   U2727 : OAI21_X1 port map( B1 => n2995, B2 => n2996, A => n2946, ZN => n2963
                           );
   U2728 : NOR3_X1 port map( A1 => n2972, A2 => n2989, A3 => n2983, ZN => n2946
                           );
   U2729 : INV_X1 port map( A => n2974, ZN => n2983);
   U2730 : XNOR2_X1 port map( A => n2997, B => n2998, ZN => n2974);
   U2731 : XOR2_X1 port map( A => ADD_RD1(2), B => CWP_2_port, Z => n2997);
   U2732 : INV_X1 port map( A => n2973, ZN => n2989);
   U2733 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(2), ZN => n2973);
   U2734 : XNOR2_X1 port map( A => n2999, B => n3000, ZN => n2972);
   U2735 : XOR2_X1 port map( A => n1489, B => ADD_RD1(1), Z => n3000);
   U2736 : OAI221_X1 port map( B1 => n1980, B2 => n2802, C1 => n1872, C2 => 
                           n2801, A => n3001, ZN => n2996);
   U2737 : AOI22_X1 port map( A1 => n2798, A2 => n3053, B1 => n2046, B2 => 
                           n3077, ZN => n3001);
   U2738 : NOR3_X1 port map( A1 => n3002, A2 => n3003, A3 => n3004, ZN => n2799
                           );
   U2739 : NOR3_X1 port map( A1 => n3004, A2 => n3002, A3 => n3005, ZN => n2798
                           );
   U2740 : OAI221_X1 port map( B1 => n1891, B2 => n2797, C1 => n3113, C2 => 
                           n2796, A => n3007, ZN => n2995);
   U2741 : AOI22_X1 port map( A1 => n2793, A2 => n1840, B1 => n2045, B2 => 
                           n3116, ZN => n3007);
   U2742 : NOR3_X1 port map( A1 => n3006, A2 => n3004, A3 => n3005, ZN => n2794
                           );
   U2743 : NOR3_X1 port map( A1 => n3004, A2 => n3003, A3 => n3006, ZN => n2793
                           );
   U2744 : INV_X1 port map( A => n3002, ZN => n3006);
   U2745 : XOR2_X1 port map( A => n1490, B => n2988, Z => n3004);
   U2746 : INV_X1 port map( A => n3003, ZN => n3005);
   U2747 : XNOR2_X1 port map( A => n3008, B => n3009, ZN => n3003);
   U2748 : XOR2_X1 port map( A => n1487, B => ADD_RD1(3), Z => n3009);
   U2749 : XOR2_X1 port map( A => n3010, B => n1486, Z => n3002);
   U2750 : OAI22_X1 port map( A1 => n3008, A2 => n3011, B1 => n1487, B2 => 
                           n3012, ZN => n3010);
   U2751 : AND2_X1 port map( A1 => n3011, A2 => n3008, ZN => n3012);
   U2752 : INV_X1 port map( A => ADD_RD1(3), ZN => n3011);
   U2753 : AOI21_X1 port map( B1 => n2998, B2 => ADD_RD1(2), A => n3013, ZN => 
                           n3008);
   U2754 : INV_X1 port map( A => n3014, ZN => n3013);
   U2755 : OAI21_X1 port map( B1 => ADD_RD1(2), B2 => n2998, A => CWP_2_port, 
                           ZN => n3014);
   U2756 : OAI21_X1 port map( B1 => n3015, B2 => n2990, A => n3016, ZN => n2998
                           );
   U2757 : INV_X1 port map( A => n3017, ZN => n3016);
   U2758 : AOI21_X1 port map( B1 => n3015, B2 => n2990, A => n1489, ZN => n3017
                           );
   U2759 : INV_X1 port map( A => ADD_RD1(1), ZN => n2990);
   U2760 : INV_X1 port map( A => n2999, ZN => n3015);
   U2761 : NOR2_X1 port map( A1 => n2988, A2 => n1490, ZN => n2999);
   U2762 : INV_X1 port map( A => ADD_RD1(0), ZN => n2988);
   U2763 : OAI221_X1 port map( B1 => n3018, B2 => n3019, C1 => n1266, C2 => 
                           n2115, A => n3020, ZN => U3_U22_Z_3);
   U2764 : NOR2_X1 port map( A1 => U3_U23_Z_0, A2 => n3021, ZN => n3020);
   U2765 : INV_X1 port map( A => n2141, ZN => n3021);
   U2766 : NAND4_X1 port map( A1 => n2408, A2 => ENABLE, A3 => CALL, A4 => 
                           n2155, ZN => n2141);
   U2767 : OAI21_X1 port map( B1 => n3022, B2 => n2115, A => n3023, ZN => 
                           U3_U23_Z_0);
   U2768 : NAND3_X1 port map( A1 => n2103, A2 => ENABLE, A3 => n2408, ZN => 
                           n3023);
   U2769 : AND2_X1 port map( A1 => n2154, A2 => n2144, ZN => n2103);
   U2770 : AND2_X1 port map( A1 => RET, A2 => n2143, ZN => n2154);
   U2771 : INV_X1 port map( A => FILL_port, ZN => n3022);
   U2772 : INV_X1 port map( A => n2130, ZN => n2115);
   U2773 : INV_X1 port map( A => ADD_WR(3), ZN => n3018);
   U2774 : NOR2_X1 port map( A1 => n3024, A2 => n3019, ZN => U3_U22_Z_2);
   U2775 : INV_X1 port map( A => ADD_WR(2), ZN => n3024);
   U2776 : NOR2_X1 port map( A1 => n2175, A2 => n3019, ZN => U3_U22_Z_1);
   U2777 : INV_X1 port map( A => ADD_WR(1), ZN => n2175);
   U2778 : NOR2_X1 port map( A1 => n2171, A2 => n3019, ZN => U3_U22_Z_0);
   U2779 : NAND3_X1 port map( A1 => n2408, A2 => n2180, A3 => n2409, ZN => 
                           n3019);
   U2780 : AND4_X1 port map( A1 => WR, A2 => ENABLE, A3 => n2144, A4 => n2142, 
                           ZN => n2409);
   U2781 : INV_X1 port map( A => RET, ZN => n2142);
   U2782 : NAND2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n2180);
   U2783 : INV_X1 port map( A => ADD_WR(0), ZN => n2171);
   U2784 : OAI21_X1 port map( B1 => n2130, B2 => n2133, A => n3025, ZN => N202)
                           ;
   U2785 : NAND4_X1 port map( A1 => RET, A2 => n2144, A3 => ENABLE, A4 => n3026
                           , ZN => n3025);
   U2786 : NOR2_X1 port map( A1 => n2143, A2 => n2132, ZN => n3026);
   U2787 : NAND2_X1 port map( A1 => n3281, A2 => n3282, ZN => n2143);
   U2788 : NAND2_X1 port map( A1 => FILL_port, A2 => n2093, ZN => n2133);
   U2789 : NOR2_X1 port map( A1 => n1944, A2 => n3283, ZN => FILL_port);
   U2790 : OAI33_X1 port map( A1 => n2130, A2 => RESET, A3 => n1266, B1 => 
                           n3027, B2 => n3028, B3 => n2132, ZN => N201);
   U2791 : NAND2_X1 port map( A1 => n2408, A2 => n2093, ZN => n2132);
   U2792 : INV_X1 port map( A => RESET, ZN => n2093);
   U2793 : NOR2_X1 port map( A1 => n3283, A2 => n3286, ZN => n2408);
   U2794 : INV_X1 port map( A => ENABLE, ZN => n3028);
   U2795 : OR2_X1 port map( A1 => n2144, A2 => n2155, ZN => n3027);
   U2796 : NAND2_X1 port map( A1 => n3284, A2 => n3285, ZN => n2155);
   U2797 : INV_X1 port map( A => CALL, ZN => n2144);
   U2798 : NAND2_X1 port map( A1 => n3283, A2 => n1944, ZN => n1266);
   U2799 : NOR2_X1 port map( A1 => n1889, A2 => n2111, ZN => n2130);
   U2800 : NAND2_X1 port map( A1 => n1495, A2 => n1494, ZN => n2111);

end SYN_BEHAVIORAL;


library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_959;

architecture SYN_BEHAVIORAL of FA_959 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_958;

architecture SYN_BEHAVIORAL of FA_958 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_957;

architecture SYN_BEHAVIORAL of FA_957 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : CLKBUF_X1 port map( A => n5, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_956;

architecture SYN_BEHAVIORAL of FA_956 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n7);
   U2 : AOI22_X1 port map( A1 => B, A2 => n6, B1 => Ci, B2 => n5, ZN => n4);
   U5 : INV_X1 port map( A => n4, ZN => Co);
   U6 : CLKBUF_X1 port map( A => A, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_955;

architecture SYN_BEHAVIORAL of FA_955 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : AOI21_X1 port map( B1 => Ci, B2 => n6, A => n4, ZN => n2);
   U3 : INV_X1 port map( A => n2, ZN => Co);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U5 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_954;

architecture SYN_BEHAVIORAL of FA_954 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net148237, net155753, n4, n5, n6 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => net148237, B => net155753, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net155753);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net148237);
   U5 : NOR2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U6 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U7 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_953;

architecture SYN_BEHAVIORAL of FA_953 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U3 : AOI21_X1 port map( B1 => Ci, B2 => n5, A => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_952;

architecture SYN_BEHAVIORAL of FA_952 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_951;

architecture SYN_BEHAVIORAL of FA_951 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U3 : INV_X1 port map( A => n6, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U5 : AOI21_X1 port map( B1 => Ci, B2 => n5, A => n4, ZN => n2);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_950;

architecture SYN_BEHAVIORAL of FA_950 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_949;

architecture SYN_BEHAVIORAL of FA_949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_948;

architecture SYN_BEHAVIORAL of FA_948 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_947;

architecture SYN_BEHAVIORAL of FA_947 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_946;

architecture SYN_BEHAVIORAL of FA_946 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_945;

architecture SYN_BEHAVIORAL of FA_945 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_944;

architecture SYN_BEHAVIORAL of FA_944 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_943;

architecture SYN_BEHAVIORAL of FA_943 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_942;

architecture SYN_BEHAVIORAL of FA_942 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_941;

architecture SYN_BEHAVIORAL of FA_941 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_940;

architecture SYN_BEHAVIORAL of FA_940 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_939;

architecture SYN_BEHAVIORAL of FA_939 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_938;

architecture SYN_BEHAVIORAL of FA_938 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_937;

architecture SYN_BEHAVIORAL of FA_937 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_936;

architecture SYN_BEHAVIORAL of FA_936 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_935;

architecture SYN_BEHAVIORAL of FA_935 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : INV_X1 port map( A => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_934;

architecture SYN_BEHAVIORAL of FA_934 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : INV_X1 port map( A => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_933;

architecture SYN_BEHAVIORAL of FA_933 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_932;

architecture SYN_BEHAVIORAL of FA_932 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_931;

architecture SYN_BEHAVIORAL of FA_931 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_930;

architecture SYN_BEHAVIORAL of FA_930 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_929;

architecture SYN_BEHAVIORAL of FA_929 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_928;

architecture SYN_BEHAVIORAL of FA_928 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_927;

architecture SYN_BEHAVIORAL of FA_927 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_926;

architecture SYN_BEHAVIORAL of FA_926 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_925;

architecture SYN_BEHAVIORAL of FA_925 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_924;

architecture SYN_BEHAVIORAL of FA_924 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : INV_X1 port map( A => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_923;

architecture SYN_BEHAVIORAL of FA_923 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_922;

architecture SYN_BEHAVIORAL of FA_922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_921;

architecture SYN_BEHAVIORAL of FA_921 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_920;

architecture SYN_BEHAVIORAL of FA_920 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_919 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_919;

architecture SYN_BEHAVIORAL of FA_919 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_918 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_918;

architecture SYN_BEHAVIORAL of FA_918 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : BUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_917 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_917;

architecture SYN_BEHAVIORAL of FA_917 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_916 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_916;

architecture SYN_BEHAVIORAL of FA_916 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_915 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_915;

architecture SYN_BEHAVIORAL of FA_915 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_914 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_914;

architecture SYN_BEHAVIORAL of FA_914 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_913 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_913;

architecture SYN_BEHAVIORAL of FA_913 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_912 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_912;

architecture SYN_BEHAVIORAL of FA_912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_911 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_911;

architecture SYN_BEHAVIORAL of FA_911 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_910 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_910;

architecture SYN_BEHAVIORAL of FA_910 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_909 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_909;

architecture SYN_BEHAVIORAL of FA_909 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_908 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_908;

architecture SYN_BEHAVIORAL of FA_908 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_907 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_907;

architecture SYN_BEHAVIORAL of FA_907 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_906 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_906;

architecture SYN_BEHAVIORAL of FA_906 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_905 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_905;

architecture SYN_BEHAVIORAL of FA_905 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_904 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_904;

architecture SYN_BEHAVIORAL of FA_904 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_903 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_903;

architecture SYN_BEHAVIORAL of FA_903 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_902 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_902;

architecture SYN_BEHAVIORAL of FA_902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_901 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_901;

architecture SYN_BEHAVIORAL of FA_901 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_900 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_900;

architecture SYN_BEHAVIORAL of FA_900 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_899 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_899;

architecture SYN_BEHAVIORAL of FA_899 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_898 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_898;

architecture SYN_BEHAVIORAL of FA_898 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_897 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_897;

architecture SYN_BEHAVIORAL of FA_897 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_896 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_896;

architecture SYN_BEHAVIORAL of FA_896 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_895 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_895;

architecture SYN_BEHAVIORAL of FA_895 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_894 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_894;

architecture SYN_BEHAVIORAL of FA_894 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_893 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_893;

architecture SYN_BEHAVIORAL of FA_893 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_892 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_892;

architecture SYN_BEHAVIORAL of FA_892 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_891 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_891;

architecture SYN_BEHAVIORAL of FA_891 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n6, ZN => S);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U3 : AND2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : AOI21_X1 port map( B1 => n6, B2 => n7, A => n5, ZN => Co);
   U5 : INV_X1 port map( A => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n4, ZN => n9);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U8 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_890 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_890;

architecture SYN_BEHAVIORAL of FA_890 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net140187, net140208, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net140208, B => net140187, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => net140208);
   U2 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U4 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n5);
   U6 : XOR2_X1 port map( A => B, B => A, Z => net140187);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_889 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_889;

architecture SYN_BEHAVIORAL of FA_889 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_888 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_888;

architecture SYN_BEHAVIORAL of FA_888 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_887 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_887;

architecture SYN_BEHAVIORAL of FA_887 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_886 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_886;

architecture SYN_BEHAVIORAL of FA_886 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_885 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_885;

architecture SYN_BEHAVIORAL of FA_885 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_884 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_884;

architecture SYN_BEHAVIORAL of FA_884 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_883 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_883;

architecture SYN_BEHAVIORAL of FA_883 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_882 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_882;

architecture SYN_BEHAVIORAL of FA_882 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_881 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_881;

architecture SYN_BEHAVIORAL of FA_881 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_880 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_880;

architecture SYN_BEHAVIORAL of FA_880 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => n7, Z => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : OAI22_X1 port map( A1 => n5, A2 => n7, B1 => n6, B2 => n4, ZN => Co);
   U4 : INV_X1 port map( A => B, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_879 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_879;

architecture SYN_BEHAVIORAL of FA_879 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_878 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_878;

architecture SYN_BEHAVIORAL of FA_878 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => n8, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_877 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_877;

architecture SYN_BEHAVIORAL of FA_877 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U4 : INV_X32 port map( A => A, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n6);
   U6 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_876 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_876;

architecture SYN_BEHAVIORAL of FA_876 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_875 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_875;

architecture SYN_BEHAVIORAL of FA_875 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_874 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_874;

architecture SYN_BEHAVIORAL of FA_874 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_873 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_873;

architecture SYN_BEHAVIORAL of FA_873 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_872 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_872;

architecture SYN_BEHAVIORAL of FA_872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_871 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_871;

architecture SYN_BEHAVIORAL of FA_871 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_870 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_870;

architecture SYN_BEHAVIORAL of FA_870 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_869 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_869;

architecture SYN_BEHAVIORAL of FA_869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_868 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_868;

architecture SYN_BEHAVIORAL of FA_868 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_867 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_867;

architecture SYN_BEHAVIORAL of FA_867 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => n8);
   U4 : INV_X32 port map( A => A, ZN => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_866 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_866;

architecture SYN_BEHAVIORAL of FA_866 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_865 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_865;

architecture SYN_BEHAVIORAL of FA_865 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_864 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_864;

architecture SYN_BEHAVIORAL of FA_864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_863 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_863;

architecture SYN_BEHAVIORAL of FA_863 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_862 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_862;

architecture SYN_BEHAVIORAL of FA_862 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_861 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_861;

architecture SYN_BEHAVIORAL of FA_861 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_860 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_860;

architecture SYN_BEHAVIORAL of FA_860 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_859 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_859;

architecture SYN_BEHAVIORAL of FA_859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_858 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_858;

architecture SYN_BEHAVIORAL of FA_858 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_857 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_857;

architecture SYN_BEHAVIORAL of FA_857 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_856 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_856;

architecture SYN_BEHAVIORAL of FA_856 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_855 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_855;

architecture SYN_BEHAVIORAL of FA_855 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_854 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_854;

architecture SYN_BEHAVIORAL of FA_854 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U4 : INV_X32 port map( A => A, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_853 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_853;

architecture SYN_BEHAVIORAL of FA_853 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_852 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_852;

architecture SYN_BEHAVIORAL of FA_852 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_851 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_851;

architecture SYN_BEHAVIORAL of FA_851 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_850 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_850;

architecture SYN_BEHAVIORAL of FA_850 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_849 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_849;

architecture SYN_BEHAVIORAL of FA_849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_848 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_848;

architecture SYN_BEHAVIORAL of FA_848 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_847 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_847;

architecture SYN_BEHAVIORAL of FA_847 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_846 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_846;

architecture SYN_BEHAVIORAL of FA_846 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_845 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_845;

architecture SYN_BEHAVIORAL of FA_845 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_844 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_844;

architecture SYN_BEHAVIORAL of FA_844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_843 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_843;

architecture SYN_BEHAVIORAL of FA_843 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_842 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_842;

architecture SYN_BEHAVIORAL of FA_842 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_841 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_841;

architecture SYN_BEHAVIORAL of FA_841 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_840 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_840;

architecture SYN_BEHAVIORAL of FA_840 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_839 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_839;

architecture SYN_BEHAVIORAL of FA_839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_838 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_838;

architecture SYN_BEHAVIORAL of FA_838 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_837 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_837;

architecture SYN_BEHAVIORAL of FA_837 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_836 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_836;

architecture SYN_BEHAVIORAL of FA_836 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_835 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_835;

architecture SYN_BEHAVIORAL of FA_835 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_834 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_834;

architecture SYN_BEHAVIORAL of FA_834 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_833 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_833;

architecture SYN_BEHAVIORAL of FA_833 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_832 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_832;

architecture SYN_BEHAVIORAL of FA_832 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_831 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_831;

architecture SYN_BEHAVIORAL of FA_831 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_830 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_830;

architecture SYN_BEHAVIORAL of FA_830 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_829 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_829;

architecture SYN_BEHAVIORAL of FA_829 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_828 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_828;

architecture SYN_BEHAVIORAL of FA_828 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_827 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_827;

architecture SYN_BEHAVIORAL of FA_827 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_826 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_826;

architecture SYN_BEHAVIORAL of FA_826 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_825 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_825;

architecture SYN_BEHAVIORAL of FA_825 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_824 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_824;

architecture SYN_BEHAVIORAL of FA_824 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n10, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n10, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : CLKBUF_X1 port map( A => Ci, Z => n7);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_823 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_823;

architecture SYN_BEHAVIORAL of FA_823 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_822 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_822;

architecture SYN_BEHAVIORAL of FA_822 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_821 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_821;

architecture SYN_BEHAVIORAL of FA_821 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_820 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_820;

architecture SYN_BEHAVIORAL of FA_820 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_819 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_819;

architecture SYN_BEHAVIORAL of FA_819 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_818 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_818;

architecture SYN_BEHAVIORAL of FA_818 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XOR2_X1 port map( A => B, B => n8, Z => n4);
   U3 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n7, B2 => n4, ZN => Co);
   U5 : INV_X1 port map( A => n5, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_817 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_817;

architecture SYN_BEHAVIORAL of FA_817 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_816 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_816;

architecture SYN_BEHAVIORAL of FA_816 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_815 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_815;

architecture SYN_BEHAVIORAL of FA_815 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_814 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_814;

architecture SYN_BEHAVIORAL of FA_814 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_813 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_813;

architecture SYN_BEHAVIORAL of FA_813 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_812 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_812;

architecture SYN_BEHAVIORAL of FA_812 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_811 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_811;

architecture SYN_BEHAVIORAL of FA_811 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_810 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_810;

architecture SYN_BEHAVIORAL of FA_810 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_809 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_809;

architecture SYN_BEHAVIORAL of FA_809 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_808 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_808;

architecture SYN_BEHAVIORAL of FA_808 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_807 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_807;

architecture SYN_BEHAVIORAL of FA_807 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_806 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_806;

architecture SYN_BEHAVIORAL of FA_806 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_805 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_805;

architecture SYN_BEHAVIORAL of FA_805 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_804 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_804;

architecture SYN_BEHAVIORAL of FA_804 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_803 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_803;

architecture SYN_BEHAVIORAL of FA_803 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_802 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_802;

architecture SYN_BEHAVIORAL of FA_802 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_801 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_801;

architecture SYN_BEHAVIORAL of FA_801 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_800 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_800;

architecture SYN_BEHAVIORAL of FA_800 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_799 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_799;

architecture SYN_BEHAVIORAL of FA_799 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_798 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_798;

architecture SYN_BEHAVIORAL of FA_798 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_797 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_797;

architecture SYN_BEHAVIORAL of FA_797 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_796 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_796;

architecture SYN_BEHAVIORAL of FA_796 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_795 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_795;

architecture SYN_BEHAVIORAL of FA_795 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_794 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_794;

architecture SYN_BEHAVIORAL of FA_794 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_793 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_793;

architecture SYN_BEHAVIORAL of FA_793 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_792 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_792;

architecture SYN_BEHAVIORAL of FA_792 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_791 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_791;

architecture SYN_BEHAVIORAL of FA_791 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_790 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_790;

architecture SYN_BEHAVIORAL of FA_790 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_789 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_789;

architecture SYN_BEHAVIORAL of FA_789 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U4 : INV_X32 port map( A => A, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_788 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_788;

architecture SYN_BEHAVIORAL of FA_788 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_787 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_787;

architecture SYN_BEHAVIORAL of FA_787 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_786 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_786;

architecture SYN_BEHAVIORAL of FA_786 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_785 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_785;

architecture SYN_BEHAVIORAL of FA_785 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_784 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_784;

architecture SYN_BEHAVIORAL of FA_784 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_783 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_783;

architecture SYN_BEHAVIORAL of FA_783 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_782 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_782;

architecture SYN_BEHAVIORAL of FA_782 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_781 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_781;

architecture SYN_BEHAVIORAL of FA_781 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_780 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_780;

architecture SYN_BEHAVIORAL of FA_780 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_779 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_779;

architecture SYN_BEHAVIORAL of FA_779 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_778 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_778;

architecture SYN_BEHAVIORAL of FA_778 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_777 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_777;

architecture SYN_BEHAVIORAL of FA_777 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_776 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_776;

architecture SYN_BEHAVIORAL of FA_776 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_775 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_775;

architecture SYN_BEHAVIORAL of FA_775 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_774 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_774;

architecture SYN_BEHAVIORAL of FA_774 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_773 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_773;

architecture SYN_BEHAVIORAL of FA_773 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_772 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_772;

architecture SYN_BEHAVIORAL of FA_772 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_771 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_771;

architecture SYN_BEHAVIORAL of FA_771 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_770 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_770;

architecture SYN_BEHAVIORAL of FA_770 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_769 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_769;

architecture SYN_BEHAVIORAL of FA_769 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : CLKBUF_X1 port map( A => n8, Z => n5);
   U4 : INV_X1 port map( A => n9, ZN => Co);
   U5 : INV_X1 port map( A => A, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_768 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_768;

architecture SYN_BEHAVIORAL of FA_768 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_767 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_767;

architecture SYN_BEHAVIORAL of FA_767 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_766 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_766;

architecture SYN_BEHAVIORAL of FA_766 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_765 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_765;

architecture SYN_BEHAVIORAL of FA_765 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_764 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_764;

architecture SYN_BEHAVIORAL of FA_764 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_763 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_763;

architecture SYN_BEHAVIORAL of FA_763 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_762 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_762;

architecture SYN_BEHAVIORAL of FA_762 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_761 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_761;

architecture SYN_BEHAVIORAL of FA_761 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_760 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_760;

architecture SYN_BEHAVIORAL of FA_760 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_759 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_759;

architecture SYN_BEHAVIORAL of FA_759 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_758 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_758;

architecture SYN_BEHAVIORAL of FA_758 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_757 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_757;

architecture SYN_BEHAVIORAL of FA_757 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_756 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_756;

architecture SYN_BEHAVIORAL of FA_756 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_755 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_755;

architecture SYN_BEHAVIORAL of FA_755 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_754 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_754;

architecture SYN_BEHAVIORAL of FA_754 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_753 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_753;

architecture SYN_BEHAVIORAL of FA_753 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_752 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_752;

architecture SYN_BEHAVIORAL of FA_752 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_751 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_751;

architecture SYN_BEHAVIORAL of FA_751 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_750 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_750;

architecture SYN_BEHAVIORAL of FA_750 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_749 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_749;

architecture SYN_BEHAVIORAL of FA_749 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_748 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_748;

architecture SYN_BEHAVIORAL of FA_748 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_747 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_747;

architecture SYN_BEHAVIORAL of FA_747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_746 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_746;

architecture SYN_BEHAVIORAL of FA_746 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_745 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_745;

architecture SYN_BEHAVIORAL of FA_745 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_744 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_744;

architecture SYN_BEHAVIORAL of FA_744 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_743 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_743;

architecture SYN_BEHAVIORAL of FA_743 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_742 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_742;

architecture SYN_BEHAVIORAL of FA_742 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_741 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_741;

architecture SYN_BEHAVIORAL of FA_741 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_740 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_740;

architecture SYN_BEHAVIORAL of FA_740 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_739 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_739;

architecture SYN_BEHAVIORAL of FA_739 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_738 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_738;

architecture SYN_BEHAVIORAL of FA_738 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_737 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_737;

architecture SYN_BEHAVIORAL of FA_737 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_736 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_736;

architecture SYN_BEHAVIORAL of FA_736 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_735 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_735;

architecture SYN_BEHAVIORAL of FA_735 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_734 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_734;

architecture SYN_BEHAVIORAL of FA_734 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_733 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_733;

architecture SYN_BEHAVIORAL of FA_733 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_732 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_732;

architecture SYN_BEHAVIORAL of FA_732 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_731 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_731;

architecture SYN_BEHAVIORAL of FA_731 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_730 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_730;

architecture SYN_BEHAVIORAL of FA_730 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_729 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_729;

architecture SYN_BEHAVIORAL of FA_729 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_728 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_728;

architecture SYN_BEHAVIORAL of FA_728 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_727 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_727;

architecture SYN_BEHAVIORAL of FA_727 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_726 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_726;

architecture SYN_BEHAVIORAL of FA_726 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_725 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_725;

architecture SYN_BEHAVIORAL of FA_725 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_724 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_724;

architecture SYN_BEHAVIORAL of FA_724 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_723 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_723;

architecture SYN_BEHAVIORAL of FA_723 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_722 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_722;

architecture SYN_BEHAVIORAL of FA_722 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_721 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_721;

architecture SYN_BEHAVIORAL of FA_721 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_720 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_720;

architecture SYN_BEHAVIORAL of FA_720 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_719 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_719;

architecture SYN_BEHAVIORAL of FA_719 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_718 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_718;

architecture SYN_BEHAVIORAL of FA_718 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_717 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_717;

architecture SYN_BEHAVIORAL of FA_717 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_716 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_716;

architecture SYN_BEHAVIORAL of FA_716 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_715 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_715;

architecture SYN_BEHAVIORAL of FA_715 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_714 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_714;

architecture SYN_BEHAVIORAL of FA_714 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_713 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_713;

architecture SYN_BEHAVIORAL of FA_713 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_712 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_712;

architecture SYN_BEHAVIORAL of FA_712 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_711 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_711;

architecture SYN_BEHAVIORAL of FA_711 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_710 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_710;

architecture SYN_BEHAVIORAL of FA_710 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_709 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_709;

architecture SYN_BEHAVIORAL of FA_709 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_708 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_708;

architecture SYN_BEHAVIORAL of FA_708 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_707 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_707;

architecture SYN_BEHAVIORAL of FA_707 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n8, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_706 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_706;

architecture SYN_BEHAVIORAL of FA_706 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n9);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n8, A2 => Ci, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_705 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_705;

architecture SYN_BEHAVIORAL of FA_705 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_704 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_704;

architecture SYN_BEHAVIORAL of FA_704 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_703 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_703;

architecture SYN_BEHAVIORAL of FA_703 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_702 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_702;

architecture SYN_BEHAVIORAL of FA_702 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_701 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_701;

architecture SYN_BEHAVIORAL of FA_701 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_700 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_700;

architecture SYN_BEHAVIORAL of FA_700 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_699 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_699;

architecture SYN_BEHAVIORAL of FA_699 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_698 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_698;

architecture SYN_BEHAVIORAL of FA_698 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_697 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_697;

architecture SYN_BEHAVIORAL of FA_697 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_696 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_696;

architecture SYN_BEHAVIORAL of FA_696 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_695 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_695;

architecture SYN_BEHAVIORAL of FA_695 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_694 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_694;

architecture SYN_BEHAVIORAL of FA_694 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_693 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_693;

architecture SYN_BEHAVIORAL of FA_693 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n10, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : CLKBUF_X1 port map( A => n10, Z => n7);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_692 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_692;

architecture SYN_BEHAVIORAL of FA_692 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_691 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_691;

architecture SYN_BEHAVIORAL of FA_691 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_690 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_690;

architecture SYN_BEHAVIORAL of FA_690 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_689 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_689;

architecture SYN_BEHAVIORAL of FA_689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_688 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_688;

architecture SYN_BEHAVIORAL of FA_688 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_687 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_687;

architecture SYN_BEHAVIORAL of FA_687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_686 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_686;

architecture SYN_BEHAVIORAL of FA_686 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_685 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_685;

architecture SYN_BEHAVIORAL of FA_685 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_684 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_684;

architecture SYN_BEHAVIORAL of FA_684 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_683 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_683;

architecture SYN_BEHAVIORAL of FA_683 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_682 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_682;

architecture SYN_BEHAVIORAL of FA_682 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_681 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_681;

architecture SYN_BEHAVIORAL of FA_681 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_680 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_680;

architecture SYN_BEHAVIORAL of FA_680 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_679 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_679;

architecture SYN_BEHAVIORAL of FA_679 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_678 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_678;

architecture SYN_BEHAVIORAL of FA_678 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_677 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_677;

architecture SYN_BEHAVIORAL of FA_677 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_676 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_676;

architecture SYN_BEHAVIORAL of FA_676 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_675 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_675;

architecture SYN_BEHAVIORAL of FA_675 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_674 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_674;

architecture SYN_BEHAVIORAL of FA_674 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_673 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_673;

architecture SYN_BEHAVIORAL of FA_673 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_672 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_672;

architecture SYN_BEHAVIORAL of FA_672 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_671 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_671;

architecture SYN_BEHAVIORAL of FA_671 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_670 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_670;

architecture SYN_BEHAVIORAL of FA_670 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_669 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_669;

architecture SYN_BEHAVIORAL of FA_669 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_668 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_668;

architecture SYN_BEHAVIORAL of FA_668 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_667 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_667;

architecture SYN_BEHAVIORAL of FA_667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_666 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_666;

architecture SYN_BEHAVIORAL of FA_666 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_665 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_665;

architecture SYN_BEHAVIORAL of FA_665 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_664 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_664;

architecture SYN_BEHAVIORAL of FA_664 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_663 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_663;

architecture SYN_BEHAVIORAL of FA_663 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_662 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_662;

architecture SYN_BEHAVIORAL of FA_662 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_661 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_661;

architecture SYN_BEHAVIORAL of FA_661 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_660 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_660;

architecture SYN_BEHAVIORAL of FA_660 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_659 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_659;

architecture SYN_BEHAVIORAL of FA_659 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_658 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_658;

architecture SYN_BEHAVIORAL of FA_658 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_657 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_657;

architecture SYN_BEHAVIORAL of FA_657 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_656 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_656;

architecture SYN_BEHAVIORAL of FA_656 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_655 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_655;

architecture SYN_BEHAVIORAL of FA_655 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_654 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_654;

architecture SYN_BEHAVIORAL of FA_654 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_653 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_653;

architecture SYN_BEHAVIORAL of FA_653 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_652 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_652;

architecture SYN_BEHAVIORAL of FA_652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_651 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_651;

architecture SYN_BEHAVIORAL of FA_651 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_650 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_650;

architecture SYN_BEHAVIORAL of FA_650 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_649 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_649;

architecture SYN_BEHAVIORAL of FA_649 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : OAI22_X1 port map( A1 => n5, A2 => n7, B1 => n6, B2 => n4, ZN => Co);
   U4 : INV_X1 port map( A => B, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_648 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_648;

architecture SYN_BEHAVIORAL of FA_648 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_647 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_647;

architecture SYN_BEHAVIORAL of FA_647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_646 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_646;

architecture SYN_BEHAVIORAL of FA_646 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_645 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_645;

architecture SYN_BEHAVIORAL of FA_645 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U1 : XOR2_X1 port map( A => B, B => n8, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n4, B2 => n7, ZN => Co);
   U5 : INV_X1 port map( A => n5, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_644 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_644;

architecture SYN_BEHAVIORAL of FA_644 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_643 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_643;

architecture SYN_BEHAVIORAL of FA_643 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_642 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_642;

architecture SYN_BEHAVIORAL of FA_642 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_641 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_641;

architecture SYN_BEHAVIORAL of FA_641 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_640 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_640;

architecture SYN_BEHAVIORAL of FA_640 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_639 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_639;

architecture SYN_BEHAVIORAL of FA_639 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_638 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_638;

architecture SYN_BEHAVIORAL of FA_638 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_637 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_637;

architecture SYN_BEHAVIORAL of FA_637 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_636 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_636;

architecture SYN_BEHAVIORAL of FA_636 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_635 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_635;

architecture SYN_BEHAVIORAL of FA_635 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_634 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_634;

architecture SYN_BEHAVIORAL of FA_634 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_633 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_633;

architecture SYN_BEHAVIORAL of FA_633 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_632 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_632;

architecture SYN_BEHAVIORAL of FA_632 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_631 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_631;

architecture SYN_BEHAVIORAL of FA_631 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_630 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_630;

architecture SYN_BEHAVIORAL of FA_630 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_629 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_629;

architecture SYN_BEHAVIORAL of FA_629 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_628 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_628;

architecture SYN_BEHAVIORAL of FA_628 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_627 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_627;

architecture SYN_BEHAVIORAL of FA_627 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_626 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_626;

architecture SYN_BEHAVIORAL of FA_626 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_625 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_625;

architecture SYN_BEHAVIORAL of FA_625 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_624 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_624;

architecture SYN_BEHAVIORAL of FA_624 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_623 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_623;

architecture SYN_BEHAVIORAL of FA_623 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_622 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_622;

architecture SYN_BEHAVIORAL of FA_622 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_621 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_621;

architecture SYN_BEHAVIORAL of FA_621 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_620 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_620;

architecture SYN_BEHAVIORAL of FA_620 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_619 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_619;

architecture SYN_BEHAVIORAL of FA_619 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U2 : INV_X32 port map( A => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n8);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : AOI22_X1 port map( A1 => n9, A2 => A, B1 => Ci, B2 => n7, ZN => n6);
   U6 : INV_X1 port map( A => n6, ZN => Co);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_618 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_618;

architecture SYN_BEHAVIORAL of FA_618 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_617 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_617;

architecture SYN_BEHAVIORAL of FA_617 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_616 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_616;

architecture SYN_BEHAVIORAL of FA_616 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_615 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_615;

architecture SYN_BEHAVIORAL of FA_615 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_614 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_614;

architecture SYN_BEHAVIORAL of FA_614 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_613 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_613;

architecture SYN_BEHAVIORAL of FA_613 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_612 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_612;

architecture SYN_BEHAVIORAL of FA_612 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_611 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_611;

architecture SYN_BEHAVIORAL of FA_611 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_610 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_610;

architecture SYN_BEHAVIORAL of FA_610 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_609 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_609;

architecture SYN_BEHAVIORAL of FA_609 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_608 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_608;

architecture SYN_BEHAVIORAL of FA_608 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n8);
   U2 : OR2_X1 port map( A1 => n10, A2 => n4, ZN => n6);
   U4 : INV_X1 port map( A => A, ZN => n10);
   U5 : INV_X1 port map( A => n8, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U7 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n7);
   U8 : XNOR2_X1 port map( A => B, B => n10, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => n8, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_538;

architecture SYN_BEHAVIORAL of FA_538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_537;

architecture SYN_BEHAVIORAL of FA_537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => n8, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => n8, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n8, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n9, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n9);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : CLKBUF_X1 port map( A => Ci, Z => n7);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U8 : INV_X1 port map( A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n7, A2 => n9, B1 => n8, B2 => n5, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => B, B => n9, Z => n4);
   U4 : XOR2_X1 port map( A => B, B => n9, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n6, ZN => n7);
   U7 : INV_X1 port map( A => Ci, ZN => n8);
   U8 : INV_X1 port map( A => A, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n12, n13 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n12, A2 => n5, ZN => n6);
   U2 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => S);
   U4 : INV_X1 port map( A => n12, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n10);
   U7 : CLKBUF_X1 port map( A => n12, Z => n8);
   U8 : CLKBUF_X1 port map( A => B, Z => n9);
   U9 : XNOR2_X1 port map( A => B, B => n10, ZN => n12);
   U10 : INV_X1 port map( A => n13, ZN => Co);
   U11 : AOI22_X1 port map( A1 => n9, A2 => A, B1 => n8, B2 => Ci, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n8, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n11, n12, n13 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n11, A2 => n5, ZN => n6);
   U2 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => S);
   U4 : INV_X1 port map( A => n11, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n13);
   U7 : NAND2_X1 port map( A1 => n12, A2 => A, ZN => n8);
   U8 : NAND2_X1 port map( A1 => n11, A2 => Ci, ZN => n9);
   U9 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => Co);
   U10 : XNOR2_X1 port map( A => B, B => n13, ZN => n11);
   U11 : CLKBUF_X1 port map( A => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n13, n14 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => n11, Z => n4);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n13, ZN => n6);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => S);
   U5 : INV_X1 port map( A => Ci, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n11);
   U7 : CLKBUF_X1 port map( A => Ci, Z => n8);
   U8 : CLKBUF_X1 port map( A => B, Z => n9);
   U9 : CLKBUF_X1 port map( A => n13, Z => n10);
   U10 : XNOR2_X1 port map( A => B, B => n11, ZN => n13);
   U11 : INV_X1 port map( A => n14, ZN => Co);
   U12 : AOI22_X1 port map( A1 => n9, A2 => A, B1 => n10, B2 => n8, ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U2 : INV_X32 port map( A => n11, ZN => n4);
   U3 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => n11, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n11);
   U6 : NAND2_X1 port map( A1 => n10, A2 => A, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n6, A2 => Ci, ZN => n8);
   U8 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Co);
   U9 : CLKBUF_X1 port map( A => B, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : CLKBUF_X1 port map( A => n9, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n9);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => n4, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n8, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : XOR2_X1 port map( A => B, B => n9, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n9, B1 => n7, B2 => n4, ZN => Co);
   U5 : INV_X1 port map( A => n5, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n9);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n8, B2 => n4, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);
   U6 : CLKBUF_X1 port map( A => n5, Z => n8);
   U7 : CLKBUF_X1 port map( A => B, Z => n6);
   U8 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n9, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net145650, net145834, net145860, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U2 : AND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U3 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net145860);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U6 : CLKBUF_X1 port map( A => n6, Z => net145834);
   U7 : CLKBUF_X1 port map( A => B, Z => n7);
   U8 : INV_X1 port map( A => net145860, ZN => net145650);
   U9 : NOR2_X1 port map( A1 => net145650, A2 => net145834, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n8);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => n6, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n9, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => n9, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n9);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U1 : CLKBUF_X1 port map( A => n10, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U4 : INV_X1 port map( A => A, ZN => n9);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n10, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net144039, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : NOR2_X1 port map( A1 => n4, A2 => Ci, ZN => n6);
   U3 : XNOR2_X1 port map( A => net144039, B => Ci, ZN => S);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net144039);
   U6 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136396, net145762, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : BUF_X1 port map( A => Ci, Z => net136396);
   U3 : XNOR2_X1 port map( A => net145762, B => net136396, ZN => S);
   U4 : OR2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => n7, A => n5, ZN => n6);
   U6 : INV_X1 port map( A => n6, ZN => Co);
   U7 : AND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U8 : XNOR2_X1 port map( A => n4, B => A, ZN => net145762);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net158915, net158910, n4, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : OR2_X1 port map( A1 => n9, A2 => n6, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => n8, ZN => n6);
   U4 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);
   U5 : INV_X1 port map( A => n4, ZN => net158910);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U7 : CLKBUF_X1 port map( A => n7, Z => net158915);
   U8 : CLKBUF_X1 port map( A => B, Z => n8);
   U9 : NOR2_X1 port map( A1 => net158915, A2 => net158910, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_14;

architecture SYN_STRUCTURAL of RCA_NBIT64_14 is

   component FA_833
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_834
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_835
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_836
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_837
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_838
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_839
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_840
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_841
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_842
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_843
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_844
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_845
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_846
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_847
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_848
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_849
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_850
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_851
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_852
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_853
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_854
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_855
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_856
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_857
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_858
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_859
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_860
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_861
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_862
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_863
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_864
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_865
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_866
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_867
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_868
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_869
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_870
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_871
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_872
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_873
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_874
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_875
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_876
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_877
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_878
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_879
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_880
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_881
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_882
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_883
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_884
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_885
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_886
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_887
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_888
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_889
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_890
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_891
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_892
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_893
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_894
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_895
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_896
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_896 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_895 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_894 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_893 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_892 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_891 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_890 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_889 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_888 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_887 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_886 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_885 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_884 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_883 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_882 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_881 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_880 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_879 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_878 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_877 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_876 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_875 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_874 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_873 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_872 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_871 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_870 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_869 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_868 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_867 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_866 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_865 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_864 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_863 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_862 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_861 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_860 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_859 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_858 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_857 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_856 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_855 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_854 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_853 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_852 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_851 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_850 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_849 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_848 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_847 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_846 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_845 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_844 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_843 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_842 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_841 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_840 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_839 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_838 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_837 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_836 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_835 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_834 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_833 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_13;

architecture SYN_STRUCTURAL of RCA_NBIT64_13 is

   component FA_769
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_770
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_771
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_772
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_773
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_774
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_775
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_776
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_777
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_778
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_779
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_780
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_781
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_782
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_783
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_784
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_785
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_786
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_787
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_788
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_789
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_790
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_791
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_792
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_793
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_794
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_795
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_796
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_797
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_798
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_799
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_800
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_801
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_802
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_803
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_804
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_805
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_806
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_807
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_808
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_809
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_810
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_811
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_812
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_813
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_814
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_815
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_816
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_817
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_818
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_819
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_820
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_821
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_822
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_823
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_824
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_825
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_826
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_827
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_828
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_829
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_830
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_831
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_832
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_832 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_831 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_830 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_829 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_828 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_827 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_826 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_825 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_824 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_823 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_822 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_821 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_820 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_819 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_818 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_817 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_816 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_815 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_814 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_813 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_812 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_811 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_810 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_809 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_808 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_807 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_806 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_805 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_804 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_803 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_802 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_801 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_800 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_799 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_798 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_797 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_796 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_795 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_794 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_793 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_792 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_791 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_790 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_789 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_788 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_787 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_786 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_785 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_784 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_783 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_782 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_781 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_780 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_779 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_778 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_777 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_776 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_775 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_774 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_773 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_772 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_771 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_770 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_769 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_12;

architecture SYN_STRUCTURAL of RCA_NBIT64_12 is

   component FA_705
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_706
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_707
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_708
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_709
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_710
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_711
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_712
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_713
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_714
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_715
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_716
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_717
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_718
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_719
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_720
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_721
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_722
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_723
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_724
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_725
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_726
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_727
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_728
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_729
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_730
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_731
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_732
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_733
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_734
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_735
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_736
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_737
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_738
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_739
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_740
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_741
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_742
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_743
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_744
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_745
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_746
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_747
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_748
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_749
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_750
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_751
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_752
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_753
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_754
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_755
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_756
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_757
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_758
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_759
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_760
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_761
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_762
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_763
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_764
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_765
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_766
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_767
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_768
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_768 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_767 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_766 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_765 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_764 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_763 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_762 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_761 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_760 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_759 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_758 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_757 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_756 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_755 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_754 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_753 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_752 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_751 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_750 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_749 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_748 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_747 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_746 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_745 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_744 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_743 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_742 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_741 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_740 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_739 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_738 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_737 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_736 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_735 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_734 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_733 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_732 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_731 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_730 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_729 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_728 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_727 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_726 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_725 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_724 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_723 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_722 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_721 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_720 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_719 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_718 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_717 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_716 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_715 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_714 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_713 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_712 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_711 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_710 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_709 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_708 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_707 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_706 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_705 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_11;

architecture SYN_STRUCTURAL of RCA_NBIT64_11 is

   component FA_641
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_642
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_643
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_644
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_645
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_646
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_647
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_648
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_649
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_650
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_651
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_652
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_653
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_654
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_655
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_656
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_657
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_658
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_659
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_660
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_661
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_662
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_663
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_664
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_665
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_666
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_667
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_668
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_669
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_670
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_671
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_672
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_673
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_674
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_675
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_676
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_677
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_678
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_679
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_680
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_681
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_682
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_683
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_684
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_685
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_686
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_687
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_688
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_689
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_690
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_691
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_692
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_693
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_694
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_695
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_696
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_697
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_698
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_699
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_700
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_701
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_702
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_703
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_704
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_704 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_703 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_702 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_701 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_700 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_699 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_698 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_697 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_696 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_695 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_694 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_693 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_692 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_691 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_690 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_689 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_688 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_687 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_686 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_685 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_684 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_683 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_682 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_681 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_680 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_679 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_678 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_677 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_676 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_675 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_674 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_673 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_672 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_671 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_670 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_669 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_668 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_667 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_666 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_665 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_664 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_663 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_662 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_661 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_660 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_659 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_658 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_657 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_656 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_655 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_654 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_653 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_652 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_651 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_650 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_649 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_648 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_647 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_646 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_645 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_644 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_643 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_642 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_641 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_10;

architecture SYN_STRUCTURAL of RCA_NBIT64_10 is

   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_608
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_609
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_610
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_611
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_612
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_613
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_614
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_615
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_616
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_617
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_618
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_619
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_620
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_621
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_622
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_623
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_624
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_625
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_626
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_627
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_628
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_629
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_630
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_631
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_632
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_633
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_634
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_635
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_636
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_637
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_638
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_639
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_640
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_640 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_639 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_638 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_637 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_636 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_635 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_634 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_633 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_632 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_631 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_630 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_629 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_628 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_627 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_626 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_625 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_624 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_623 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_622 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_621 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_620 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_619 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_618 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_617 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_616 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_615 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_614 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_613 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_612 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_611 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_610 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_609 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_608 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_607 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_606 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_605 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_604 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_603 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_602 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_601 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_600 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_599 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_598 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_597 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_596 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_595 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_594 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_593 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_592 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_591 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_590 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_589 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_588 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_587 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_586 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_585 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_584 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_583 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_582 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_581 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_580 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_579 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_578 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_577 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_9;

architecture SYN_STRUCTURAL of RCA_NBIT64_9 is

   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_576 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_575 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_574 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_573 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_572 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_571 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_570 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_569 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_568 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_567 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_566 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_565 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_564 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_563 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_562 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_561 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_560 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_559 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_558 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_557 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_556 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_555 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_554 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_553 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_552 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_551 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_550 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_549 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_548 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_547 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_546 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_545 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_544 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_543 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_542 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_541 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_540 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_539 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_538 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_537 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_536 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_535 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_534 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_533 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_532 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_531 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_530 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_529 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_528 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_527 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_526 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_525 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_524 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_523 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_522 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_521 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_520 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_519 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_518 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_517 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_516 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_515 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_514 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_513 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_8;

architecture SYN_STRUCTURAL of RCA_NBIT64_8 is

   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_512 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_511 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_510 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_509 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_508 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_507 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_506 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_505 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_504 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_503 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_502 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_501 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_500 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_499 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_498 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_497 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_496 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_495 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_494 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_493 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_492 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_491 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_490 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_489 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_488 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_487 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_486 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_485 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_484 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_483 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_482 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_481 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_480 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_479 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_478 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_477 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_476 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_475 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_474 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_473 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_472 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_471 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_470 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_469 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_468 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_467 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_466 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_465 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_464 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_463 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_462 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_461 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_460 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_459 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_458 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_457 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_456 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_455 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_454 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_453 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_452 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_451 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_450 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_449 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_7;

architecture SYN_STRUCTURAL of RCA_NBIT64_7 is

   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_448 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_447 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_446 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_445 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_444 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_443 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_442 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_441 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_440 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_439 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_438 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_437 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_436 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_435 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_434 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_433 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_432 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_431 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_430 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_429 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_428 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_427 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_426 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_425 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_424 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_423 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_422 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_421 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_420 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_419 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_418 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_417 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_416 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_415 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_414 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_413 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_412 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_411 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_410 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_409 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_408 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_407 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_406 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_405 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_404 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_403 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_402 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_401 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_400 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_399 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_398 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_397 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_396 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_395 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_394 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_393 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_392 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_391 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_390 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_389 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_388 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_387 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_386 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_385 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_6;

architecture SYN_STRUCTURAL of RCA_NBIT64_6 is

   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_384 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_383 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_382 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_381 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_380 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_379 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_378 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_377 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_376 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_375 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_374 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_373 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_372 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_371 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_370 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_369 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_368 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_367 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_366 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_365 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_364 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_363 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_362 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_361 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_360 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_359 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_358 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_357 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_356 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_355 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_354 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_353 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_352 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_351 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_350 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_349 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_348 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_347 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_346 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_345 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_344 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_343 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_342 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_341 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_340 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_339 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_338 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_337 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_336 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_335 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_334 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_333 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_332 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_331 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_330 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_329 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_328 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_327 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_326 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_325 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_324 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_323 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_322 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_321 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_5;

architecture SYN_STRUCTURAL of RCA_NBIT64_5 is

   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_320 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_319 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_318 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_317 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_316 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_315 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_314 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_313 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_312 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_311 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_310 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_309 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_308 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_307 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_306 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_305 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_304 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_303 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_302 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_301 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_300 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_299 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_298 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_297 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_296 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_295 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_294 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_293 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_292 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_291 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_290 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_289 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_288 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_287 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_286 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_285 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_284 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_283 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_282 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_281 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_280 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_279 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_278 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_277 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_276 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_275 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_274 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_273 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_272 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_271 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_270 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_269 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_268 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_267 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_266 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_265 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_264 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_263 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_262 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_261 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_260 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_259 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_258 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_257 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_4;

architecture SYN_STRUCTURAL of RCA_NBIT64_4 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_256 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_255 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_254 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_253 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_252 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_251 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_250 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_249 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_248 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_247 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_246 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_245 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_244 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_243 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_242 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_241 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_240 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_239 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_238 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_237 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_236 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_235 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_234 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_233 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_232 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_231 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_230 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_229 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_228 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_227 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_226 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_225 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_224 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_223 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_222 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_221 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_220 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_219 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_218 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_217 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_216 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_215 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_214 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_213 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_212 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_211 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_210 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_209 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_208 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_207 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_206 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_205 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_204 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_203 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_202 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_201 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_200 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_199 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_198 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_197 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_196 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_195 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_194 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_193 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_3;

architecture SYN_STRUCTURAL of RCA_NBIT64_3 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_192 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_191 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_190 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_189 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_188 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_187 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_186 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_185 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_184 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_183 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_182 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_181 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_180 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_179 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_178 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_177 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_176 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_175 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_174 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_173 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_172 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_171 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_170 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_169 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_168 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_167 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_166 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_165 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_164 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_163 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_162 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_161 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_160 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_159 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_158 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_157 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_156 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_155 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_154 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_153 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_152 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_151 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_150 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_149 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_148 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_147 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_146 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_145 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_144 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_143 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_142 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_141 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_140 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_139 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_138 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_137 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_136 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_135 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_134 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_133 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_132 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_131 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_130 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_129 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_2;

architecture SYN_STRUCTURAL of RCA_NBIT64_2 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_124 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_123 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_122 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_121 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_120 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_119 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_118 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_117 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_116 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_115 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_114 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_113 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_112 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_111 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_110 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_109 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_108 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_107 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_106 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_105 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_104 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_103 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_102 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_101 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_100 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_99 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_98 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_97 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_96 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_95 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_94 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_93 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_92 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_91 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_90 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_89 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_88 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_87 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_86 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_85 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_84 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_83 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_82 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_81 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_80 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_79 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_78 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_77 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_76 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_75 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_74 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_73 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_72 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_71 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_70 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_69 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_68 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_67 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_66 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_65 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_1;

architecture SYN_STRUCTURAL of RCA_NBIT64_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_60 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_59 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_58 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_57 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => CTMP_8_port);
   FAI_9 : FA_56 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8), 
                           Co => CTMP_9_port);
   FAI_10 : FA_55 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9),
                           Co => CTMP_10_port);
   FAI_11 : FA_54 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_53 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_52 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_51 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_50 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_49 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_48 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_47 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_46 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_45 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_44 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_43 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_42 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_41 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_40 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_39 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_38 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_37 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_36 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_35 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_34 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_33 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_32 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_31 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_30 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_29 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_28 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_27 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_26 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_25 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_24 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_23 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_22 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_21 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_20 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_19 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_18 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_17 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_16 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_15 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_14 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_13 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_12 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_11 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_10 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_9 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_8 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_7 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_6 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_5 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_4 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_3 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_2 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_15 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_15;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n13, n23, n67, n88, net129597, net129596, net129594, net129593, 
      net129630, net129629, net129700, net129703, net129717, net129720, 
      net129973, net129993, net129991, net129985, net129983, net132879, 
      net136168, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => net136168, Z => n138);
   U2 : BUF_X1 port map( A => net129703, Z => net129720);
   U3 : CLKBUF_X1 port map( A => n178, Z => n186);
   U4 : BUF_X2 port map( A => n178, Z => n185);
   U5 : CLKBUF_X1 port map( A => n178, Z => n184);
   U6 : BUF_X4 port map( A => n183, Z => n181);
   U7 : BUF_X2 port map( A => sel(2), Z => n183);
   U8 : CLKBUF_X1 port map( A => net132879, Z => n139);
   U9 : INV_X1 port map( A => A1(8), ZN => n155);
   U10 : NOR2_X1 port map( A1 => n157, A2 => n171, ZN => n149);
   U11 : INV_X1 port map( A => A3(8), ZN => n157);
   U12 : NOR2_X1 port map( A1 => n162, A2 => n140, ZN => n150);
   U13 : INV_X1 port map( A => A1(5), ZN => n162);
   U14 : NOR2_X1 port map( A1 => n163, A2 => n171, ZN => n151);
   U15 : INV_X1 port map( A => A3(5), ZN => n163);
   U16 : NAND2_X1 port map( A1 => A3(6), A2 => n144, ZN => n169);
   U17 : INV_X1 port map( A => A1(6), ZN => n164);
   U18 : INV_X1 port map( A => A3(2), ZN => n165);
   U19 : INV_X1 port map( A => A1(3), ZN => n159);
   U20 : NOR3_X1 port map( A1 => n137, A2 => n148, A3 => n149, ZN => n9);
   U21 : NOR2_X1 port map( A1 => n155, A2 => n140, ZN => n148);
   U22 : NOR3_X1 port map( A1 => n136, A2 => n150, A3 => n151, ZN => n23);
   U23 : NOR2_X1 port map( A1 => n172, A2 => n147, ZN => n13);
   U24 : OAI21_X1 port map( B1 => n164, B2 => n140, A => n169, ZN => n147);
   U25 : BUF_X1 port map( A => net129596, Z => net129991);
   U26 : BUF_X1 port map( A => n174, Z => net129973);
   U27 : AND2_X1 port map( A1 => A2(5), A2 => net129703, ZN => n136);
   U28 : AND2_X1 port map( A1 => A2(8), A2 => net129594, ZN => n137);
   U29 : AND2_X2 port map( A1 => n138, A2 => n139, ZN => n144);
   U30 : NOR2_X1 port map( A1 => n170, A2 => n165, ZN => n166);
   U31 : CLKBUF_X1 port map( A => n156, Z => n140);
   U32 : INV_X1 port map( A => n160, ZN => n141);
   U33 : BUF_X1 port map( A => net129703, Z => net129593);
   U34 : CLKBUF_X1 port map( A => n139, Z => n142);
   U35 : INV_X1 port map( A => n140, ZN => n143);
   U36 : NOR2_X1 port map( A1 => n159, A2 => n156, ZN => n145);
   U37 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => O(2));
   U38 : AOI21_X1 port map( B1 => A1(2), B2 => net129629, A => n167, ZN => n152
                           );
   U39 : INV_X1 port map( A => n88, ZN => n167);
   U40 : NOR2_X1 port map( A1 => n146, A2 => n145, ZN => n67);
   U41 : INV_X1 port map( A => n158, ZN => n173);
   U42 : CLKBUF_X1 port map( A => net129703, Z => net129594);
   U43 : BUF_X1 port map( A => net129593, Z => net129596);
   U44 : BUF_X1 port map( A => net129594, Z => net129597);
   U45 : CLKBUF_X1 port map( A => net129596, Z => net129993);
   U46 : CLKBUF_X1 port map( A => net129993, Z => net129983);
   U47 : BUF_X4 port map( A => net129991, Z => net129985);
   U48 : CLKBUF_X1 port map( A => net129629, Z => net129630);
   U49 : BUF_X4 port map( A => n143, Z => net129700);
   U50 : OR2_X1 port map( A1 => sel(1), A2 => n154, ZN => n156);
   U51 : AOI21_X1 port map( B1 => A2(2), B2 => n141, A => n166, ZN => n153);
   U52 : NAND3_X1 port map( A1 => net132879, A2 => net136168, A3 => A3(3), ZN 
                           => n168);
   U53 : INV_X1 port map( A => n156, ZN => net129629);
   U54 : CLKBUF_X1 port map( A => n175, Z => net129717);
   U55 : NAND2_X1 port map( A1 => net136168, A2 => net132879, ZN => n158);
   U56 : INV_X1 port map( A => n173, ZN => n170);
   U57 : INV_X1 port map( A => n173, ZN => n171);
   U58 : INV_X1 port map( A => n158, ZN => n177);
   U59 : INV_X1 port map( A => n140, ZN => n175);
   U60 : INV_X1 port map( A => sel(0), ZN => n154);
   U61 : INV_X1 port map( A => n154, ZN => net132879);
   U62 : CLKBUF_X1 port map( A => net129700, Z => n176);
   U63 : INV_X2 port map( A => n170, ZN => n174);
   U64 : BUF_X1 port map( A => sel(1), Z => net136168);
   U65 : INV_X1 port map( A => A2(3), ZN => n161);
   U66 : NAND2_X1 port map( A1 => n154, A2 => sel(1), ZN => n160);
   U67 : INV_X1 port map( A => n160, ZN => net129703);
   U68 : OAI21_X1 port map( B1 => n160, B2 => n161, A => n168, ZN => n146);
   U69 : AND2_X1 port map( A1 => A2(6), A2 => net129720, ZN => n172);
   U70 : BUF_X2 port map( A => n183, Z => n180);
   U71 : NOR3_X1 port map( A1 => n138, A2 => n182, A3 => n142, ZN => n178);
   U72 : BUF_X1 port map( A => n184, Z => n187);
   U73 : NAND2_X1 port map( A1 => n309, A2 => n308, ZN => O(9));
   U74 : AOI22_X1 port map( A1 => A0(9), A2 => n185, B1 => n182, B2 => A4(9), 
                           ZN => n309);
   U75 : AOI22_X1 port map( A1 => A0(4), A2 => n184, B1 => A4(4), B2 => n180, 
                           ZN => n274);
   U76 : AOI22_X1 port map( A1 => A0(5), A2 => n187, B1 => A4(5), B2 => n181, 
                           ZN => n295);
   U77 : NAND2_X1 port map( A1 => n304, A2 => n13, ZN => O(6));
   U78 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(10));
   U79 : AOI22_X1 port map( A1 => A0(10), A2 => n184, B1 => A4(10), B2 => n181,
                           ZN => n191);
   U80 : AOI22_X1 port map( A1 => A0(7), A2 => n185, B1 => A4(7), B2 => n181, 
                           ZN => n306);
   U81 : AOI22_X1 port map( A1 => A0(8), A2 => n185, B1 => A4(8), B2 => n181, 
                           ZN => n307);
   U82 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(13));
   U83 : AOI22_X1 port map( A1 => A0(13), A2 => n184, B1 => A4(13), B2 => n181,
                           ZN => n197);
   U84 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(11));
   U85 : AOI22_X1 port map( A1 => A0(11), A2 => n184, B1 => A4(11), B2 => n181,
                           ZN => n193);
   U86 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(21));
   U87 : AOI22_X1 port map( A1 => A0(21), A2 => n185, B1 => A4(21), B2 => n181,
                           ZN => n215);
   U88 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(14));
   U89 : AOI22_X1 port map( A1 => A0(14), A2 => n184, B1 => A4(14), B2 => n181,
                           ZN => n199);
   U90 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(20));
   U91 : AOI22_X1 port map( A1 => A0(20), A2 => n185, B1 => A4(20), B2 => n181,
                           ZN => n213);
   U92 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(22));
   U93 : AOI22_X1 port map( A1 => A0(22), A2 => n185, B1 => A4(22), B2 => n181,
                           ZN => n217);
   U94 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(15));
   U95 : AOI22_X1 port map( A1 => A0(15), A2 => n184, B1 => A4(15), B2 => n181,
                           ZN => n201);
   U96 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(19));
   U97 : AOI22_X1 port map( A1 => A0(19), A2 => n184, B1 => A4(19), B2 => n181,
                           ZN => n209);
   U98 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(12));
   U99 : AOI22_X1 port map( A1 => A0(12), A2 => n184, B1 => A4(12), B2 => n181,
                           ZN => n195);
   U100 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(18));
   U101 : AOI22_X1 port map( A1 => A0(18), A2 => n184, B1 => A4(18), B2 => n181
                           , ZN => n207);
   U102 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(23));
   U103 : AOI22_X1 port map( A1 => A0(23), A2 => n185, B1 => A4(23), B2 => n181
                           , ZN => n219);
   U104 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(16));
   U105 : AOI22_X1 port map( A1 => A0(16), A2 => n184, B1 => A4(16), B2 => n181
                           , ZN => n203);
   U106 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(17));
   U107 : AOI22_X1 port map( A1 => A0(17), A2 => n184, B1 => A4(17), B2 => n181
                           , ZN => n205);
   U108 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(24));
   U109 : AOI22_X1 port map( A1 => A0(24), A2 => n185, B1 => A4(24), B2 => n181
                           , ZN => n221);
   U110 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(34));
   U111 : AOI22_X1 port map( A1 => A0(34), A2 => n186, B1 => A4(34), B2 => n180
                           , ZN => n241);
   U112 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(25));
   U113 : AOI22_X1 port map( A1 => A0(25), A2 => n185, B1 => A4(25), B2 => n181
                           , ZN => n223);
   U114 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(26));
   U115 : AOI22_X1 port map( A1 => A0(26), A2 => n185, B1 => A4(26), B2 => n181
                           , ZN => n225);
   U116 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(27));
   U117 : AOI22_X1 port map( A1 => A0(27), A2 => n185, B1 => A4(27), B2 => n181
                           , ZN => n227);
   U118 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(35));
   U119 : AOI22_X1 port map( A1 => A0(35), A2 => n186, B1 => A4(35), B2 => n180
                           , ZN => n243);
   U120 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(28));
   U121 : AOI22_X1 port map( A1 => A0(28), A2 => n185, B1 => A4(28), B2 => n181
                           , ZN => n229);
   U122 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(29));
   U123 : AOI22_X1 port map( A1 => A0(29), A2 => n185, B1 => A4(29), B2 => n181
                           , ZN => n231);
   U124 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(36));
   U125 : AOI22_X1 port map( A1 => A0(36), A2 => n186, B1 => A4(36), B2 => n180
                           , ZN => n245);
   U126 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(30));
   U127 : AOI22_X1 port map( A1 => A0(30), A2 => n185, B1 => A4(30), B2 => n181
                           , ZN => n233);
   U128 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(31));
   U129 : AOI22_X1 port map( A1 => A0(31), A2 => n186, B1 => A4(31), B2 => n181
                           , ZN => n235);
   U130 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(37));
   U131 : AOI22_X1 port map( A1 => A0(37), A2 => n186, B1 => A4(37), B2 => n179
                           , ZN => n247);
   U132 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(32));
   U133 : AOI22_X1 port map( A1 => A0(32), A2 => n186, B1 => A4(32), B2 => n181
                           , ZN => n237);
   U134 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(33));
   U135 : AOI22_X1 port map( A1 => A0(33), A2 => n186, B1 => A4(33), B2 => n181
                           , ZN => n239);
   U136 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(38));
   U137 : AOI22_X1 port map( A1 => A0(38), A2 => n186, B1 => A4(38), B2 => n179
                           , ZN => n249);
   U138 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(39));
   U139 : AOI22_X1 port map( A1 => A0(39), A2 => n186, B1 => A4(39), B2 => n179
                           , ZN => n251);
   U140 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => O(40));
   U141 : AOI22_X1 port map( A1 => A0(40), A2 => n186, B1 => A4(40), B2 => n179
                           , ZN => n254);
   U142 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => O(41));
   U143 : AOI22_X1 port map( A1 => A0(41), A2 => n186, B1 => A4(41), B2 => n179
                           , ZN => n256);
   U144 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => O(42));
   U145 : AOI22_X1 port map( A1 => A0(42), A2 => n185, B1 => A4(42), B2 => n179
                           , ZN => n258);
   U146 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => O(43));
   U147 : AOI22_X1 port map( A1 => A0(43), A2 => n186, B1 => A4(43), B2 => n179
                           , ZN => n260);
   U148 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => O(44));
   U149 : AOI22_X1 port map( A1 => A0(44), A2 => n185, B1 => A4(44), B2 => n180
                           , ZN => n262);
   U150 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => O(45));
   U151 : AOI22_X1 port map( A1 => A0(45), A2 => n186, B1 => A4(45), B2 => n180
                           , ZN => n264);
   U152 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => O(46));
   U153 : AOI22_X1 port map( A1 => A0(46), A2 => n185, B1 => A4(46), B2 => n180
                           , ZN => n266);
   U154 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => O(47));
   U155 : AOI22_X1 port map( A1 => A0(47), A2 => n186, B1 => A4(47), B2 => n180
                           , ZN => n268);
   U156 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => O(48));
   U157 : AOI22_X1 port map( A1 => A0(48), A2 => n185, B1 => A4(48), B2 => n180
                           , ZN => n270);
   U158 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => O(49));
   U159 : AOI22_X1 port map( A1 => A0(49), A2 => n186, B1 => A4(49), B2 => n180
                           , ZN => n272);
   U160 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => O(50));
   U161 : AOI22_X1 port map( A1 => A0(50), A2 => n185, B1 => A4(50), B2 => n180
                           , ZN => n276);
   U162 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => O(51));
   U163 : AOI22_X1 port map( A1 => A0(51), A2 => n186, B1 => A4(51), B2 => n179
                           , ZN => n278);
   U164 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => O(52));
   U165 : AOI22_X1 port map( A1 => A0(52), A2 => n185, B1 => A4(52), B2 => n179
                           , ZN => n280);
   U166 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => O(53));
   U167 : AOI22_X1 port map( A1 => A0(53), A2 => n187, B1 => A4(53), B2 => n179
                           , ZN => n282);
   U168 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => O(54));
   U169 : AOI22_X1 port map( A1 => A0(54), A2 => n187, B1 => A4(54), B2 => n179
                           , ZN => n284);
   U170 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => O(55));
   U171 : AOI22_X1 port map( A1 => A0(55), A2 => n187, B1 => A4(55), B2 => n179
                           , ZN => n286);
   U172 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => O(56));
   U173 : AOI22_X1 port map( A1 => A0(56), A2 => n187, B1 => A4(56), B2 => n179
                           , ZN => n288);
   U174 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => O(57));
   U175 : AOI22_X1 port map( A1 => A0(57), A2 => n187, B1 => A4(57), B2 => n179
                           , ZN => n290);
   U176 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => O(58));
   U177 : AOI22_X1 port map( A1 => A0(58), A2 => n187, B1 => A4(58), B2 => n179
                           , ZN => n292);
   U178 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => O(59));
   U179 : AOI22_X1 port map( A1 => A0(59), A2 => n187, B1 => A4(59), B2 => n180
                           , ZN => n294);
   U180 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(60));
   U181 : AOI22_X1 port map( A1 => A0(60), A2 => n187, B1 => A4(60), B2 => n179
                           , ZN => n297);
   U182 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(61));
   U183 : AOI22_X1 port map( A1 => A0(61), A2 => n187, B1 => A4(61), B2 => n179
                           , ZN => n299);
   U184 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(62));
   U185 : AOI22_X1 port map( A1 => A0(62), A2 => n187, B1 => A4(62), B2 => n179
                           , ZN => n301);
   U186 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(63));
   U187 : AOI22_X1 port map( A1 => A0(63), A2 => n187, B1 => A4(63), B2 => n179
                           , ZN => n303);
   U188 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(0));
   U189 : AOI22_X1 port map( A1 => A0(0), A2 => n184, B1 => A4(0), B2 => n179, 
                           ZN => n189);
   U190 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(1));
   U191 : AOI22_X1 port map( A1 => A0(1), A2 => n184, B1 => A4(1), B2 => n179, 
                           ZN => n211);
   U192 : AOI222_X1 port map( A1 => A1(1), A2 => n176, B1 => A3(1), B2 => n174,
                           C1 => A2(1), C2 => net129985, ZN => n210);
   U193 : CLKBUF_X1 port map( A => n181, Z => n179);
   U194 : BUF_X1 port map( A => n183, Z => n182);
   U195 : AOI222_X1 port map( A1 => A1(61), A2 => n176, B1 => A3(61), B2 => 
                           n174, C1 => A2(61), C2 => net129985, ZN => n298);
   U196 : AOI222_X1 port map( A1 => A1(58), A2 => n176, B1 => A3(58), B2 => 
                           n174, C1 => A2(58), C2 => net129985, ZN => n291);
   U197 : AOI222_X1 port map( A1 => A1(55), A2 => n176, B1 => A3(55), B2 => 
                           n144, C1 => A2(55), C2 => net129985, ZN => n285);
   U198 : AOI222_X1 port map( A1 => A1(52), A2 => n176, B1 => A3(52), B2 => 
                           n174, C1 => A2(52), C2 => net129985, ZN => n279);
   U199 : AOI222_X1 port map( A1 => A1(49), A2 => n176, B1 => A3(49), B2 => 
                           n174, C1 => A2(49), C2 => net129985, ZN => n271);
   U200 : AOI222_X1 port map( A1 => A1(46), A2 => n176, B1 => A3(46), B2 => 
                           n173, C1 => A2(46), C2 => net129985, ZN => n265);
   U201 : AOI222_X1 port map( A1 => A1(43), A2 => n176, B1 => A3(43), B2 => 
                           n174, C1 => A2(43), C2 => net129985, ZN => n259);
   U202 : AOI222_X1 port map( A1 => A1(40), A2 => n176, B1 => A3(40), B2 => 
                           n174, C1 => A2(40), C2 => net129985, ZN => n253);
   U203 : AOI222_X1 port map( A1 => A1(37), A2 => n176, B1 => A3(37), B2 => 
                           n174, C1 => A2(37), C2 => net129985, ZN => n246);
   U204 : AOI222_X1 port map( A1 => A1(34), A2 => n176, B1 => A3(34), B2 => 
                           n173, C1 => A2(34), C2 => net129985, ZN => n240);
   U205 : AOI222_X1 port map( A1 => A1(31), A2 => net129700, B1 => A3(31), B2 
                           => n144, C1 => A2(31), C2 => net129985, ZN => n234);
   U206 : AOI222_X1 port map( A1 => A1(28), A2 => net129700, B1 => A3(28), B2 
                           => n173, C1 => A2(28), C2 => net129985, ZN => n228);
   U207 : AOI222_X1 port map( A1 => A1(25), A2 => net129700, B1 => A3(25), B2 
                           => n174, C1 => A2(25), C2 => net129985, ZN => n222);
   U208 : AOI222_X1 port map( A1 => A1(22), A2 => net129700, B1 => A3(22), B2 
                           => n174, C1 => A2(22), C2 => net129985, ZN => n216);
   U209 : AOI222_X1 port map( A1 => A1(19), A2 => net129700, B1 => A3(19), B2 
                           => n144, C1 => A2(19), C2 => net129985, ZN => n208);
   U210 : AOI222_X1 port map( A1 => A1(16), A2 => net129700, B1 => A3(16), B2 
                           => net129973, C1 => A2(16), C2 => net129985, ZN => 
                           n202);
   U211 : AOI222_X1 port map( A1 => A1(13), A2 => net129700, B1 => A3(13), B2 
                           => net129973, C1 => A2(13), C2 => net129991, ZN => 
                           n196);
   U212 : AOI222_X1 port map( A1 => A1(10), A2 => net129700, B1 => A3(10), B2 
                           => n144, C1 => A2(10), C2 => net129597, ZN => n190);
   U213 : AOI222_X1 port map( A1 => A1(0), A2 => net129717, B1 => A3(0), B2 => 
                           n174, C1 => A2(0), C2 => net129985, ZN => n188);
   U214 : AOI222_X1 port map( A1 => A1(63), A2 => net129717, B1 => A3(63), B2 
                           => n144, C1 => A2(63), C2 => net129985, ZN => n302);
   U215 : AOI222_X1 port map( A1 => A1(59), A2 => net129717, B1 => A3(59), B2 
                           => n174, C1 => A2(59), C2 => net129985, ZN => n293);
   U216 : AOI222_X1 port map( A1 => A1(56), A2 => net129717, B1 => A3(56), B2 
                           => n173, C1 => A2(56), C2 => net129985, ZN => n287);
   U217 : AOI222_X1 port map( A1 => A1(53), A2 => net129717, B1 => A3(53), B2 
                           => n174, C1 => A2(53), C2 => net129985, ZN => n281);
   U218 : AOI222_X1 port map( A1 => A1(50), A2 => net129717, B1 => A3(50), B2 
                           => n144, C1 => A2(50), C2 => net129985, ZN => n275);
   U219 : AOI222_X1 port map( A1 => A1(47), A2 => net129717, B1 => A3(47), B2 
                           => n174, C1 => A2(47), C2 => net129985, ZN => n267);
   U220 : AOI222_X1 port map( A1 => A1(44), A2 => net129717, B1 => A3(44), B2 
                           => n174, C1 => A2(44), C2 => net129985, ZN => n261);
   U221 : AOI222_X1 port map( A1 => A1(41), A2 => net129717, B1 => A3(41), B2 
                           => n144, C1 => A2(41), C2 => net129985, ZN => n255);
   U222 : AOI222_X1 port map( A1 => A1(38), A2 => net129717, B1 => A3(38), B2 
                           => n144, C1 => A2(38), C2 => net129985, ZN => n248);
   U223 : AOI222_X1 port map( A1 => A1(35), A2 => net129717, B1 => A3(35), B2 
                           => n174, C1 => A2(35), C2 => net129985, ZN => n242);
   U224 : AOI222_X1 port map( A1 => A1(32), A2 => net129717, B1 => A3(32), B2 
                           => n173, C1 => A2(32), C2 => net129985, ZN => n236);
   U225 : AOI222_X1 port map( A1 => A1(29), A2 => net129717, B1 => A3(29), B2 
                           => n174, C1 => A2(29), C2 => net129985, ZN => n230);
   U226 : AOI222_X1 port map( A1 => A1(26), A2 => n175, B1 => A3(26), B2 => 
                           n173, C1 => A2(26), C2 => net129985, ZN => n224);
   U227 : AOI222_X1 port map( A1 => A1(23), A2 => net129717, B1 => A3(23), B2 
                           => n174, C1 => A2(23), C2 => net129985, ZN => n218);
   U228 : AOI222_X1 port map( A1 => A1(20), A2 => net129717, B1 => A3(20), B2 
                           => n173, C1 => A2(20), C2 => net129985, ZN => n212);
   U229 : AOI222_X1 port map( A1 => A1(17), A2 => n175, B1 => A3(17), B2 => 
                           n174, C1 => A2(17), C2 => net129985, ZN => n204);
   U230 : AOI222_X1 port map( A1 => A1(14), A2 => n175, B1 => A3(14), B2 => 
                           net129973, C1 => A2(14), C2 => net129983, ZN => n198
                           );
   U231 : AOI222_X1 port map( A1 => A1(11), A2 => n175, B1 => A3(11), B2 => 
                           n174, C1 => A2(11), C2 => net129596, ZN => n192);
   U232 : AOI222_X1 port map( A1 => A1(62), A2 => net129700, B1 => A3(62), B2 
                           => n174, C1 => A2(62), C2 => net129985, ZN => n300);
   U233 : AOI222_X1 port map( A1 => A1(60), A2 => net129700, B1 => A3(60), B2 
                           => n144, C1 => A2(60), C2 => net129985, ZN => n296);
   U234 : AOI222_X1 port map( A1 => A1(57), A2 => net129700, B1 => A3(57), B2 
                           => n174, C1 => A2(57), C2 => net129985, ZN => n289);
   U235 : AOI222_X1 port map( A1 => A1(54), A2 => net129700, B1 => A3(54), B2 
                           => n174, C1 => A2(54), C2 => net129985, ZN => n283);
   U236 : AOI222_X1 port map( A1 => A1(51), A2 => net129700, B1 => A3(51), B2 
                           => n173, C1 => A2(51), C2 => net129985, ZN => n277);
   U237 : AOI222_X1 port map( A1 => A1(48), A2 => net129700, B1 => A3(48), B2 
                           => n174, C1 => A2(48), C2 => net129985, ZN => n269);
   U238 : AOI222_X1 port map( A1 => A1(45), A2 => net129700, B1 => A3(45), B2 
                           => n174, C1 => A2(45), C2 => net129985, ZN => n263);
   U239 : AOI222_X1 port map( A1 => A1(42), A2 => net129700, B1 => A3(42), B2 
                           => n174, C1 => A2(42), C2 => net129985, ZN => n257);
   U240 : AOI222_X1 port map( A1 => A1(39), A2 => net129700, B1 => A3(39), B2 
                           => n173, C1 => A2(39), C2 => net129985, ZN => n250);
   U241 : AOI222_X1 port map( A1 => A1(36), A2 => net129700, B1 => A3(36), B2 
                           => n174, C1 => A2(36), C2 => net129985, ZN => n244);
   U242 : AOI222_X1 port map( A1 => A1(33), A2 => net129700, B1 => A3(33), B2 
                           => n174, C1 => A2(33), C2 => net129985, ZN => n238);
   U243 : AOI222_X1 port map( A1 => A1(30), A2 => net129700, B1 => A3(30), B2 
                           => n174, C1 => A2(30), C2 => net129985, ZN => n232);
   U244 : AOI222_X1 port map( A1 => A1(27), A2 => net129700, B1 => A3(27), B2 
                           => n174, C1 => A2(27), C2 => net129985, ZN => n226);
   U245 : AOI222_X1 port map( A1 => A1(24), A2 => net129700, B1 => A3(24), B2 
                           => n144, C1 => A2(24), C2 => net129985, ZN => n220);
   U246 : AOI222_X1 port map( A1 => A1(21), A2 => net129700, B1 => A3(21), B2 
                           => n173, C1 => A2(21), C2 => net129985, ZN => n214);
   U247 : AOI222_X1 port map( A1 => A1(18), A2 => net129700, B1 => A3(18), B2 
                           => n144, C1 => A2(18), C2 => net129985, ZN => n206);
   U248 : AOI222_X1 port map( A1 => A1(15), A2 => net129700, B1 => A3(15), B2 
                           => net129973, C1 => A2(15), C2 => net129983, ZN => 
                           n200);
   U249 : AOI222_X1 port map( A1 => A1(12), A2 => net129700, B1 => A3(12), B2 
                           => net129973, C1 => A2(12), C2 => net129993, ZN => 
                           n194);
   U250 : AOI222_X1 port map( A1 => A1(4), A2 => net129630, B1 => n177, B2 => 
                           A3(4), C1 => A2(4), C2 => n141, ZN => n273);
   U251 : AOI22_X1 port map( A1 => A0(6), A2 => n186, B1 => A4(6), B2 => n182, 
                           ZN => n304);
   U252 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => O(7));
   U253 : AOI222_X1 port map( A1 => A1(9), A2 => net129700, B1 => A3(9), B2 => 
                           n173, C1 => A2(9), C2 => net129593, ZN => n308);
   U254 : NAND2_X1 port map( A1 => n307, A2 => n9, ZN => O(8));
   U255 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => O(4));
   U256 : AOI222_X1 port map( A1 => A1(7), A2 => net129700, B1 => A3(7), B2 => 
                           n144, C1 => A2(7), C2 => net129720, ZN => n305);
   U257 : NAND2_X1 port map( A1 => n295, A2 => n23, ZN => O(5));
   U258 : NAND2_X1 port map( A1 => n252, A2 => n67, ZN => O(3));
   U259 : AOI22_X1 port map( A1 => A0(3), A2 => n186, B1 => A4(3), B2 => n182, 
                           ZN => n252);
   U260 : AOI22_X1 port map( A1 => A0(2), A2 => n185, B1 => A4(2), B2 => n182, 
                           ZN => n88);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_14 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_14;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_14 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => O(39));
   U2 : CLKBUF_X1 port map( A => n178, Z => n175);
   U3 : CLKBUF_X1 port map( A => n162, Z => n159);
   U4 : CLKBUF_X1 port map( A => n136, Z => n155);
   U5 : CLKBUF_X1 port map( A => n138, Z => n163);
   U6 : CLKBUF_X1 port map( A => n137, Z => n171);
   U7 : CLKBUF_X1 port map( A => n179, Z => n174);
   U8 : CLKBUF_X1 port map( A => n179, Z => n173);
   U9 : BUF_X1 port map( A => n136, Z => n154);
   U10 : BUF_X1 port map( A => n137, Z => n170);
   U11 : BUF_X1 port map( A => n138, Z => n162);
   U12 : BUF_X1 port map( A => n307, Z => n147);
   U13 : AND2_X1 port map( A1 => sel(1), A2 => n180, ZN => n136);
   U14 : NOR2_X1 port map( A1 => n180, A2 => sel(1), ZN => n137);
   U15 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U16 : BUF_X1 port map( A => sel(2), Z => n179);
   U17 : CLKBUF_X1 port map( A => sel(2), Z => n178);
   U18 : BUF_X1 port map( A => n154, Z => n152);
   U19 : BUF_X1 port map( A => n154, Z => n151);
   U20 : BUF_X1 port map( A => n162, Z => n160);
   U21 : BUF_X1 port map( A => n170, Z => n168);
   U22 : BUF_X1 port map( A => n170, Z => n167);
   U23 : BUF_X1 port map( A => n154, Z => n153);
   U24 : BUF_X1 port map( A => n162, Z => n161);
   U25 : BUF_X1 port map( A => n170, Z => n169);
   U26 : BUF_X1 port map( A => n155, Z => n148);
   U27 : BUF_X1 port map( A => n163, Z => n156);
   U28 : BUF_X1 port map( A => n171, Z => n164);
   U29 : BUF_X1 port map( A => n163, Z => n157);
   U30 : BUF_X1 port map( A => n155, Z => n149);
   U31 : BUF_X1 port map( A => n171, Z => n165);
   U32 : BUF_X1 port map( A => n163, Z => n158);
   U33 : BUF_X1 port map( A => n155, Z => n150);
   U34 : BUF_X1 port map( A => n171, Z => n166);
   U35 : BUF_X1 port map( A => n146, Z => n144);
   U36 : BUF_X1 port map( A => n147, Z => n140);
   U37 : BUF_X1 port map( A => n147, Z => n141);
   U38 : BUF_X1 port map( A => n147, Z => n142);
   U39 : BUF_X1 port map( A => n146, Z => n143);
   U40 : BUF_X1 port map( A => n146, Z => n145);
   U41 : BUF_X1 port map( A => n179, Z => n172);
   U42 : BUF_X1 port map( A => n178, Z => n177);
   U43 : BUF_X1 port map( A => n178, Z => n176);
   U44 : BUF_X1 port map( A => n307, Z => n146);
   U45 : OR3_X1 port map( A1 => sel(1), A2 => n177, A3 => sel(0), ZN => n139);
   U46 : INV_X1 port map( A => n139, ZN => n307);
   U47 : AOI22_X1 port map( A1 => A0(4), A2 => n143, B1 => A4(4), B2 => n173, 
                           ZN => n270);
   U48 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => O(6));
   U49 : AOI22_X1 port map( A1 => A0(6), A2 => n145, B1 => A4(6), B2 => n172, 
                           ZN => n302);
   U50 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161, 
                           C1 => A2(6), C2 => n153, ZN => n301);
   U51 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => O(7));
   U52 : AOI22_X1 port map( A1 => A0(7), A2 => n145, B1 => A4(7), B2 => n172, 
                           ZN => n304);
   U53 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161, 
                           C1 => A2(7), C2 => n153, ZN => n303);
   U54 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => O(8));
   U55 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161, 
                           C1 => A2(8), C2 => n153, ZN => n305);
   U56 : NAND2_X1 port map( A1 => n309, A2 => n308, ZN => O(9));
   U57 : AOI22_X1 port map( A1 => A0(9), A2 => n145, B1 => n177, B2 => A4(9), 
                           ZN => n309);
   U58 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161, 
                           C1 => A2(9), C2 => n153, ZN => n308);
   U59 : AOI22_X1 port map( A1 => A0(11), A2 => n140, B1 => A4(11), B2 => n177,
                           ZN => n186);
   U60 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => n156
                           , C1 => A2(11), C2 => n148, ZN => n185);
   U61 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => O(12));
   U62 : AOI22_X1 port map( A1 => A0(12), A2 => n140, B1 => A4(12), B2 => n176,
                           ZN => n188);
   U63 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => n156
                           , C1 => A2(12), C2 => n148, ZN => n187);
   U64 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => O(10));
   U65 : AOI22_X1 port map( A1 => A0(10), A2 => n140, B1 => A4(10), B2 => n177,
                           ZN => n184);
   U66 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => n156
                           , C1 => A2(10), C2 => n148, ZN => n183);
   U67 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => O(21));
   U68 : AOI22_X1 port map( A1 => A0(21), A2 => n141, B1 => A4(21), B2 => n176,
                           ZN => n208);
   U69 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => n157
                           , C1 => A2(21), C2 => n149, ZN => n207);
   U70 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => O(22));
   U71 : AOI22_X1 port map( A1 => A0(22), A2 => n141, B1 => A4(22), B2 => n176,
                           ZN => n210);
   U72 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => n157
                           , C1 => A2(22), C2 => n149, ZN => n209);
   U73 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => O(19));
   U74 : AOI22_X1 port map( A1 => A0(19), A2 => n140, B1 => A4(19), B2 => n176,
                           ZN => n202);
   U75 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n201);
   U76 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => O(15));
   U77 : AOI22_X1 port map( A1 => A0(15), A2 => n140, B1 => A4(15), B2 => n176,
                           ZN => n194);
   U78 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n193);
   U79 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => O(32));
   U80 : AOI22_X1 port map( A1 => A0(32), A2 => n142, B1 => A4(32), B2 => n175,
                           ZN => n232);
   U81 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => n158
                           , C1 => A2(32), C2 => n150, ZN => n231);
   U82 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => O(23));
   U83 : AOI22_X1 port map( A1 => A0(23), A2 => n141, B1 => A4(23), B2 => n175,
                           ZN => n212);
   U84 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => n157
                           , C1 => A2(23), C2 => n149, ZN => n211);
   U85 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => O(16));
   U86 : AOI22_X1 port map( A1 => A0(16), A2 => n140, B1 => A4(16), B2 => n176,
                           ZN => n196);
   U87 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n195);
   U88 : AOI22_X1 port map( A1 => A0(39), A2 => n142, B1 => A4(39), B2 => n174,
                           ZN => n246);
   U89 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => n158
                           , C1 => A2(39), C2 => n150, ZN => n245);
   U90 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => O(24));
   U91 : AOI22_X1 port map( A1 => A0(24), A2 => n141, B1 => A4(24), B2 => n175,
                           ZN => n214);
   U92 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => n157
                           , C1 => A2(24), C2 => n149, ZN => n213);
   U93 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => O(13));
   U94 : AOI22_X1 port map( A1 => A0(13), A2 => n140, B1 => A4(13), B2 => n176,
                           ZN => n190);
   U95 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => n156
                           , C1 => A2(13), C2 => n148, ZN => n189);
   U96 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => O(17));
   U97 : AOI22_X1 port map( A1 => A0(17), A2 => n140, B1 => A4(17), B2 => n176,
                           ZN => n198);
   U98 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n197);
   U99 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => O(20));
   U100 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => 
                           n157, C1 => A2(20), C2 => n149, ZN => n205);
   U101 : AOI22_X1 port map( A1 => A0(20), A2 => n141, B1 => A4(20), B2 => n176
                           , ZN => n206);
   U102 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => O(25));
   U103 : AOI22_X1 port map( A1 => A0(25), A2 => n141, B1 => A4(25), B2 => n175
                           , ZN => n216);
   U104 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => 
                           n157, C1 => A2(25), C2 => n149, ZN => n215);
   U105 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => O(14));
   U106 : AOI22_X1 port map( A1 => A0(14), A2 => n140, B1 => A4(14), B2 => n176
                           , ZN => n192);
   U107 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => 
                           n156, C1 => A2(14), C2 => n148, ZN => n191);
   U108 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => O(18));
   U109 : AOI22_X1 port map( A1 => A0(18), A2 => n140, B1 => A4(18), B2 => n176
                           , ZN => n200);
   U110 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => 
                           n156, C1 => A2(18), C2 => n148, ZN => n199);
   U111 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => O(26));
   U112 : AOI22_X1 port map( A1 => A0(26), A2 => n141, B1 => A4(26), B2 => n175
                           , ZN => n218);
   U113 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => 
                           n157, C1 => A2(26), C2 => n149, ZN => n217);
   U114 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => O(36));
   U115 : AOI22_X1 port map( A1 => A0(36), A2 => n142, B1 => A4(36), B2 => n174
                           , ZN => n240);
   U116 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n239);
   U117 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => O(27));
   U118 : AOI22_X1 port map( A1 => A0(27), A2 => n141, B1 => A4(27), B2 => n175
                           , ZN => n220);
   U119 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => 
                           n157, C1 => A2(27), C2 => n149, ZN => n219);
   U120 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => O(28));
   U121 : AOI22_X1 port map( A1 => A0(28), A2 => n141, B1 => A4(28), B2 => n175
                           , ZN => n222);
   U122 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => 
                           n157, C1 => A2(28), C2 => n149, ZN => n221);
   U123 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => O(37));
   U124 : AOI22_X1 port map( A1 => A0(37), A2 => n142, B1 => A4(37), B2 => n174
                           , ZN => n242);
   U125 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n241);
   U126 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => O(29));
   U127 : AOI22_X1 port map( A1 => A0(29), A2 => n141, B1 => A4(29), B2 => n175
                           , ZN => n224);
   U128 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => 
                           n157, C1 => A2(29), C2 => n149, ZN => n223);
   U129 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => O(30));
   U130 : AOI22_X1 port map( A1 => A0(30), A2 => n141, B1 => A4(30), B2 => n175
                           , ZN => n228);
   U131 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => 
                           n157, C1 => A2(30), C2 => n149, ZN => n227);
   U132 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => O(31));
   U133 : AOI22_X1 port map( A1 => A0(31), A2 => n142, B1 => A4(31), B2 => n175
                           , ZN => n230);
   U134 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => 
                           n158, C1 => A2(31), C2 => n150, ZN => n229);
   U135 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => O(38));
   U136 : AOI22_X1 port map( A1 => A0(38), A2 => n142, B1 => A4(38), B2 => n174
                           , ZN => n244);
   U137 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n243);
   U138 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => O(33));
   U139 : AOI22_X1 port map( A1 => A0(33), A2 => n142, B1 => A4(33), B2 => n175
                           , ZN => n234);
   U140 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => 
                           n158, C1 => A2(33), C2 => n150, ZN => n233);
   U141 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => O(34));
   U142 : AOI22_X1 port map( A1 => A0(34), A2 => n142, B1 => A4(34), B2 => n174
                           , ZN => n236);
   U143 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n235);
   U144 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => O(35));
   U145 : AOI22_X1 port map( A1 => A0(35), A2 => n142, B1 => A4(35), B2 => n174
                           , ZN => n238);
   U146 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n237);
   U147 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => O(40));
   U148 : AOI22_X1 port map( A1 => A0(40), A2 => n142, B1 => A4(40), B2 => n174
                           , ZN => n250);
   U149 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n249);
   U150 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => O(41));
   U151 : AOI22_X1 port map( A1 => A0(41), A2 => n142, B1 => A4(41), B2 => n174
                           , ZN => n252);
   U152 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n251);
   U153 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => O(42));
   U154 : AOI22_X1 port map( A1 => A0(42), A2 => n143, B1 => A4(42), B2 => n174
                           , ZN => n254);
   U155 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n253);
   U156 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => O(43));
   U157 : AOI22_X1 port map( A1 => A0(43), A2 => n143, B1 => A4(43), B2 => n174
                           , ZN => n256);
   U158 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n255);
   U159 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => O(44));
   U160 : AOI22_X1 port map( A1 => A0(44), A2 => n143, B1 => A4(44), B2 => n173
                           , ZN => n258);
   U161 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n257);
   U162 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => O(45));
   U163 : AOI22_X1 port map( A1 => A0(45), A2 => n143, B1 => A4(45), B2 => n173
                           , ZN => n260);
   U164 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n259);
   U165 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => O(46));
   U166 : AOI22_X1 port map( A1 => A0(46), A2 => n143, B1 => A4(46), B2 => n173
                           , ZN => n262);
   U167 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n261);
   U168 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => O(47));
   U169 : AOI22_X1 port map( A1 => A0(47), A2 => n143, B1 => A4(47), B2 => n173
                           , ZN => n264);
   U170 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n263);
   U171 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => O(48));
   U172 : AOI22_X1 port map( A1 => A0(48), A2 => n143, B1 => A4(48), B2 => n173
                           , ZN => n266);
   U173 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n265);
   U174 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => O(49));
   U175 : AOI22_X1 port map( A1 => A0(49), A2 => n143, B1 => A4(49), B2 => n173
                           , ZN => n268);
   U176 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n267);
   U177 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => O(50));
   U178 : AOI22_X1 port map( A1 => A0(50), A2 => n143, B1 => A4(50), B2 => n173
                           , ZN => n272);
   U179 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n271);
   U180 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => O(51));
   U181 : AOI22_X1 port map( A1 => A0(51), A2 => n143, B1 => A4(51), B2 => n173
                           , ZN => n274);
   U182 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n273);
   U183 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => O(52));
   U184 : AOI22_X1 port map( A1 => A0(52), A2 => n143, B1 => A4(52), B2 => n174
                           , ZN => n276);
   U185 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n275);
   U186 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => O(53));
   U187 : AOI22_X1 port map( A1 => A0(53), A2 => n144, B1 => A4(53), B2 => n173
                           , ZN => n278);
   U188 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n277);
   U189 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => O(54));
   U190 : AOI22_X1 port map( A1 => A0(54), A2 => n144, B1 => A4(54), B2 => n173
                           , ZN => n280);
   U191 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n279);
   U192 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => O(55));
   U193 : AOI22_X1 port map( A1 => A0(55), A2 => n144, B1 => A4(55), B2 => n173
                           , ZN => n282);
   U194 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n281);
   U195 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => O(56));
   U196 : AOI22_X1 port map( A1 => A0(56), A2 => n144, B1 => A4(56), B2 => n172
                           , ZN => n284);
   U197 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n283);
   U198 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => O(57));
   U199 : AOI22_X1 port map( A1 => A0(57), A2 => n144, B1 => A4(57), B2 => n172
                           , ZN => n286);
   U200 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n285);
   U201 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => O(58));
   U202 : AOI22_X1 port map( A1 => A0(58), A2 => n144, B1 => A4(58), B2 => n172
                           , ZN => n288);
   U203 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n287);
   U204 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => O(59));
   U205 : AOI22_X1 port map( A1 => A0(59), A2 => n144, B1 => A4(59), B2 => n172
                           , ZN => n290);
   U206 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n289);
   U207 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => O(60));
   U208 : AOI22_X1 port map( A1 => A0(60), A2 => n144, B1 => A4(60), B2 => n172
                           , ZN => n294);
   U209 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n293);
   U210 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => O(61));
   U211 : AOI22_X1 port map( A1 => A0(61), A2 => n144, B1 => A4(61), B2 => n172
                           , ZN => n296);
   U212 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n295);
   U213 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => O(62));
   U214 : AOI22_X1 port map( A1 => A0(62), A2 => n144, B1 => A4(62), B2 => n172
                           , ZN => n298);
   U215 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n297);
   U216 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => O(63));
   U217 : AOI22_X1 port map( A1 => A0(63), A2 => n144, B1 => A4(63), B2 => n172
                           , ZN => n300);
   U218 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n299);
   U219 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => O(0));
   U220 : AOI22_X1 port map( A1 => A0(0), A2 => n140, B1 => A4(0), B2 => n177, 
                           ZN => n182);
   U221 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n181);
   U222 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => O(1));
   U223 : AOI22_X1 port map( A1 => A0(1), A2 => n140, B1 => A4(1), B2 => n176, 
                           ZN => n204);
   U224 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n203);
   U225 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => O(2));
   U226 : AOI22_X1 port map( A1 => A0(2), A2 => n141, B1 => A4(2), B2 => n175, 
                           ZN => n226);
   U227 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n225);
   U228 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => O(3));
   U229 : AOI22_X1 port map( A1 => A0(3), A2 => n142, B1 => A4(3), B2 => n174, 
                           ZN => n248);
   U230 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n247);
   U231 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => O(11));
   U232 : INV_X1 port map( A => sel(0), ZN => n180);
   U233 : AOI22_X1 port map( A1 => A0(5), A2 => n144, B1 => A4(5), B2 => n172, 
                           ZN => n292);
   U234 : AOI22_X1 port map( A1 => A0(8), A2 => n145, B1 => A4(8), B2 => n172, 
                           ZN => n306);
   U235 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => O(5));
   U236 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n291);
   U237 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => O(4));
   U238 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n269);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_13 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_13;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n154, Z => n151);
   U2 : CLKBUF_X1 port map( A => n162, Z => n159);
   U3 : CLKBUF_X1 port map( A => n170, Z => n167);
   U4 : CLKBUF_X1 port map( A => n154, Z => n152);
   U5 : CLKBUF_X1 port map( A => n162, Z => n160);
   U6 : CLKBUF_X1 port map( A => n170, Z => n168);
   U7 : CLKBUF_X1 port map( A => n136, Z => n155);
   U8 : CLKBUF_X1 port map( A => n138, Z => n163);
   U9 : CLKBUF_X1 port map( A => n137, Z => n171);
   U10 : CLKBUF_X1 port map( A => n180, Z => n174);
   U11 : CLKBUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n136, Z => n154);
   U13 : BUF_X1 port map( A => n137, Z => n170);
   U14 : BUF_X1 port map( A => n138, Z => n162);
   U15 : BUF_X1 port map( A => n139, Z => n147);
   U16 : BUF_X1 port map( A => n139, Z => n146);
   U17 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U18 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n137);
   U19 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U20 : BUF_X1 port map( A => n172, Z => n180);
   U21 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n139);
   U22 : BUF_X1 port map( A => sel(2), Z => n172);
   U23 : BUF_X1 port map( A => n154, Z => n153);
   U24 : BUF_X1 port map( A => n170, Z => n169);
   U25 : BUF_X1 port map( A => n162, Z => n161);
   U26 : BUF_X1 port map( A => n171, Z => n164);
   U27 : BUF_X1 port map( A => n155, Z => n148);
   U28 : BUF_X1 port map( A => n163, Z => n156);
   U29 : BUF_X1 port map( A => n171, Z => n165);
   U30 : BUF_X1 port map( A => n163, Z => n157);
   U31 : BUF_X1 port map( A => n155, Z => n149);
   U32 : BUF_X1 port map( A => n171, Z => n166);
   U33 : BUF_X1 port map( A => n163, Z => n158);
   U34 : BUF_X1 port map( A => n155, Z => n150);
   U35 : BUF_X1 port map( A => n147, Z => n141);
   U36 : BUF_X1 port map( A => n147, Z => n142);
   U37 : BUF_X1 port map( A => n146, Z => n143);
   U38 : BUF_X1 port map( A => n146, Z => n144);
   U39 : BUF_X1 port map( A => n147, Z => n140);
   U40 : BUF_X1 port map( A => n146, Z => n145);
   U41 : BUF_X1 port map( A => n180, Z => n173);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : BUF_X1 port map( A => n179, Z => n177);
   U44 : BUF_X1 port map( A => n179, Z => n176);
   U45 : BUF_X1 port map( A => n180, Z => n175);
   U46 : AOI22_X1 port map( A1 => A0(6), A2 => n145, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U47 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161, 
                           C1 => A2(6), C2 => n153, ZN => n302);
   U48 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U49 : AOI22_X1 port map( A1 => A0(7), A2 => n145, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U50 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161, 
                           C1 => A2(7), C2 => n153, ZN => n304);
   U51 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U52 : AOI22_X1 port map( A1 => A0(8), A2 => n145, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U53 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161, 
                           C1 => A2(8), C2 => n153, ZN => n306);
   U54 : NAND2_X1 port map( A1 => n309, A2 => n308, ZN => O(9));
   U55 : AOI22_X1 port map( A1 => A0(9), A2 => n145, B1 => n178, B2 => A4(9), 
                           ZN => n309);
   U56 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161, 
                           C1 => A2(9), C2 => n153, ZN => n308);
   U57 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U58 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => n156
                           , C1 => A2(10), C2 => n148, ZN => n184);
   U59 : AOI22_X1 port map( A1 => A0(11), A2 => n140, B1 => A4(11), B2 => n178,
                           ZN => n187);
   U60 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => n156
                           , C1 => A2(11), C2 => n148, ZN => n186);
   U61 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U62 : AOI22_X1 port map( A1 => A0(12), A2 => n140, B1 => A4(12), B2 => n177,
                           ZN => n189);
   U63 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => n156
                           , C1 => A2(12), C2 => n148, ZN => n188);
   U64 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U65 : AOI22_X1 port map( A1 => A0(13), A2 => n140, B1 => A4(13), B2 => n177,
                           ZN => n191);
   U66 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => n156
                           , C1 => A2(13), C2 => n148, ZN => n190);
   U67 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U68 : AOI22_X1 port map( A1 => A0(14), A2 => n140, B1 => A4(14), B2 => n177,
                           ZN => n193);
   U69 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => n156
                           , C1 => A2(14), C2 => n148, ZN => n192);
   U70 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U71 : AOI22_X1 port map( A1 => A0(15), A2 => n140, B1 => A4(15), B2 => n177,
                           ZN => n195);
   U72 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n194);
   U73 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U74 : AOI22_X1 port map( A1 => A0(16), A2 => n140, B1 => A4(16), B2 => n177,
                           ZN => n197);
   U75 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n196);
   U76 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U77 : AOI22_X1 port map( A1 => A0(23), A2 => n141, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U78 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => n157
                           , C1 => A2(23), C2 => n149, ZN => n212);
   U79 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U80 : AOI22_X1 port map( A1 => A0(17), A2 => n140, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U81 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n198);
   U82 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U83 : AOI22_X1 port map( A1 => A0(24), A2 => n141, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U84 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => n157
                           , C1 => A2(24), C2 => n149, ZN => n214);
   U85 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U86 : AOI22_X1 port map( A1 => A0(21), A2 => n141, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U87 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => n157
                           , C1 => A2(21), C2 => n149, ZN => n208);
   U88 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U89 : AOI22_X1 port map( A1 => A0(25), A2 => n141, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U90 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => n157
                           , C1 => A2(25), C2 => n149, ZN => n216);
   U91 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U92 : AOI22_X1 port map( A1 => A0(18), A2 => n140, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U93 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => n156
                           , C1 => A2(18), C2 => n148, ZN => n200);
   U94 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U95 : AOI22_X1 port map( A1 => A0(26), A2 => n141, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U96 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => n157
                           , C1 => A2(26), C2 => n149, ZN => n218);
   U97 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U98 : AOI22_X1 port map( A1 => A0(19), A2 => n140, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U99 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n202);
   U100 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U101 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => 
                           n157, C1 => A2(22), C2 => n149, ZN => n210);
   U102 : AOI22_X1 port map( A1 => A0(22), A2 => n141, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U103 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U104 : AOI22_X1 port map( A1 => A0(27), A2 => n141, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U105 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => 
                           n157, C1 => A2(27), C2 => n149, ZN => n220);
   U106 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U107 : AOI22_X1 port map( A1 => A0(20), A2 => n141, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U108 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => 
                           n157, C1 => A2(20), C2 => n149, ZN => n206);
   U109 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U110 : AOI22_X1 port map( A1 => A0(28), A2 => n141, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U111 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => 
                           n157, C1 => A2(28), C2 => n149, ZN => n222);
   U112 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U113 : AOI22_X1 port map( A1 => A0(38), A2 => n142, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U114 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n244);
   U115 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U116 : AOI22_X1 port map( A1 => A0(29), A2 => n141, B1 => A4(29), B2 => n176
                           , ZN => n225);
   U117 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => 
                           n157, C1 => A2(29), C2 => n149, ZN => n224);
   U118 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U119 : AOI22_X1 port map( A1 => A0(30), A2 => n141, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U120 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => 
                           n157, C1 => A2(30), C2 => n149, ZN => n228);
   U121 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U122 : AOI22_X1 port map( A1 => A0(31), A2 => n142, B1 => A4(31), B2 => n176
                           , ZN => n231);
   U123 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => 
                           n158, C1 => A2(31), C2 => n150, ZN => n230);
   U124 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U125 : AOI22_X1 port map( A1 => A0(39), A2 => n142, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U126 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => 
                           n158, C1 => A2(39), C2 => n150, ZN => n246);
   U127 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U128 : AOI22_X1 port map( A1 => A0(32), A2 => n142, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U129 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => 
                           n158, C1 => A2(32), C2 => n150, ZN => n232);
   U130 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U131 : AOI22_X1 port map( A1 => A0(33), A2 => n142, B1 => A4(33), B2 => n176
                           , ZN => n235);
   U132 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => 
                           n158, C1 => A2(33), C2 => n150, ZN => n234);
   U133 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U134 : AOI22_X1 port map( A1 => A0(40), A2 => n142, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U135 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n250);
   U136 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U137 : AOI22_X1 port map( A1 => A0(34), A2 => n142, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U138 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n236);
   U139 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U140 : AOI22_X1 port map( A1 => A0(35), A2 => n142, B1 => A4(35), B2 => n175
                           , ZN => n239);
   U141 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n238);
   U142 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U143 : AOI22_X1 port map( A1 => A0(41), A2 => n142, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U144 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n252);
   U145 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U146 : AOI22_X1 port map( A1 => A0(36), A2 => n142, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U147 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n240);
   U148 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U149 : AOI22_X1 port map( A1 => A0(37), A2 => n142, B1 => A4(37), B2 => n175
                           , ZN => n243);
   U150 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n242);
   U151 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U152 : AOI22_X1 port map( A1 => A0(42), A2 => n143, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U153 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n254);
   U154 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U155 : AOI22_X1 port map( A1 => A0(43), A2 => n143, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U156 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n256);
   U157 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U158 : AOI22_X1 port map( A1 => A0(44), A2 => n143, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U159 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n258);
   U160 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U161 : AOI22_X1 port map( A1 => A0(45), A2 => n143, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U162 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n260);
   U163 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U164 : AOI22_X1 port map( A1 => A0(46), A2 => n143, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U165 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n262);
   U166 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U167 : AOI22_X1 port map( A1 => A0(47), A2 => n143, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U168 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n264);
   U169 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U170 : AOI22_X1 port map( A1 => A0(48), A2 => n143, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U171 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n266);
   U172 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U173 : AOI22_X1 port map( A1 => A0(49), A2 => n143, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U174 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n268);
   U175 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U176 : AOI22_X1 port map( A1 => A0(50), A2 => n143, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U177 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n272);
   U178 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U179 : AOI22_X1 port map( A1 => A0(51), A2 => n143, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U180 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n274);
   U181 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U182 : AOI22_X1 port map( A1 => A0(52), A2 => n143, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U183 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n276);
   U184 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U185 : AOI22_X1 port map( A1 => A0(53), A2 => n144, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U186 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n278);
   U187 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U188 : AOI22_X1 port map( A1 => A0(54), A2 => n144, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U189 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n280);
   U190 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U191 : AOI22_X1 port map( A1 => A0(55), A2 => n144, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U192 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n282);
   U193 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U194 : AOI22_X1 port map( A1 => A0(56), A2 => n144, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U195 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n284);
   U196 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U197 : AOI22_X1 port map( A1 => A0(57), A2 => n144, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U198 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n286);
   U199 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U200 : AOI22_X1 port map( A1 => A0(58), A2 => n144, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U201 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n288);
   U202 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U203 : AOI22_X1 port map( A1 => A0(63), A2 => n144, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U204 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n300);
   U205 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U206 : AOI22_X1 port map( A1 => A0(59), A2 => n144, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U207 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n290);
   U208 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U209 : AOI22_X1 port map( A1 => A0(60), A2 => n144, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U210 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n294);
   U211 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U212 : AOI22_X1 port map( A1 => A0(61), A2 => n144, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U213 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n296);
   U214 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U215 : AOI22_X1 port map( A1 => A0(62), A2 => n144, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U216 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n298);
   U217 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U218 : AOI22_X1 port map( A1 => A0(0), A2 => n140, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U219 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n182);
   U220 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U221 : AOI22_X1 port map( A1 => A0(1), A2 => n140, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U222 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n204);
   U223 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U224 : AOI22_X1 port map( A1 => A0(2), A2 => n141, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U225 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n226);
   U226 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U227 : AOI22_X1 port map( A1 => A0(3), A2 => n142, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U228 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n248);
   U229 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U230 : AOI22_X1 port map( A1 => A0(4), A2 => n143, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U231 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n270);
   U232 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U233 : AOI22_X1 port map( A1 => A0(5), A2 => n144, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U234 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n292);
   U235 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U236 : INV_X1 port map( A => sel(0), ZN => n181);
   U237 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U238 : AOI22_X1 port map( A1 => A0(10), A2 => n140, B1 => A4(10), B2 => n178
                           , ZN => n185);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_12 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_12;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n154, Z => n151);
   U2 : CLKBUF_X1 port map( A => n162, Z => n159);
   U3 : CLKBUF_X1 port map( A => n170, Z => n167);
   U4 : CLKBUF_X1 port map( A => n154, Z => n152);
   U5 : CLKBUF_X1 port map( A => n162, Z => n160);
   U6 : CLKBUF_X1 port map( A => n170, Z => n168);
   U7 : CLKBUF_X1 port map( A => n136, Z => n155);
   U8 : CLKBUF_X1 port map( A => n138, Z => n163);
   U9 : CLKBUF_X1 port map( A => n137, Z => n171);
   U10 : CLKBUF_X1 port map( A => n172, Z => n180);
   U11 : BUF_X1 port map( A => n136, Z => n154);
   U12 : BUF_X1 port map( A => n137, Z => n170);
   U13 : BUF_X1 port map( A => n138, Z => n162);
   U14 : BUF_X1 port map( A => n147, Z => n146);
   U15 : BUF_X1 port map( A => n147, Z => n145);
   U16 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U17 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n137);
   U18 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U19 : BUF_X1 port map( A => n172, Z => n179);
   U20 : BUF_X1 port map( A => sel(2), Z => n172);
   U21 : BUF_X1 port map( A => n154, Z => n153);
   U22 : BUF_X1 port map( A => n170, Z => n169);
   U23 : BUF_X1 port map( A => n162, Z => n161);
   U24 : BUF_X1 port map( A => n171, Z => n164);
   U25 : BUF_X1 port map( A => n155, Z => n148);
   U26 : BUF_X1 port map( A => n163, Z => n156);
   U27 : BUF_X1 port map( A => n171, Z => n165);
   U28 : BUF_X1 port map( A => n155, Z => n149);
   U29 : BUF_X1 port map( A => n163, Z => n157);
   U30 : BUF_X1 port map( A => n171, Z => n166);
   U31 : BUF_X1 port map( A => n155, Z => n150);
   U32 : BUF_X1 port map( A => n163, Z => n158);
   U33 : BUF_X1 port map( A => n146, Z => n140);
   U34 : BUF_X1 port map( A => n146, Z => n141);
   U35 : BUF_X1 port map( A => n145, Z => n142);
   U36 : BUF_X1 port map( A => n145, Z => n143);
   U37 : BUF_X1 port map( A => n146, Z => n139);
   U38 : BUF_X1 port map( A => n145, Z => n144);
   U39 : BUF_X1 port map( A => n179, Z => n178);
   U40 : BUF_X1 port map( A => n179, Z => n177);
   U41 : BUF_X1 port map( A => n179, Z => n176);
   U42 : BUF_X1 port map( A => n180, Z => n175);
   U43 : BUF_X1 port map( A => n180, Z => n174);
   U44 : BUF_X1 port map( A => n180, Z => n173);
   U45 : INV_X1 port map( A => sel(0), ZN => n181);
   U46 : BUF_X1 port map( A => n308, Z => n147);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U49 : AOI22_X1 port map( A1 => A0(8), A2 => n144, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U50 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161, 
                           C1 => A2(8), C2 => n153, ZN => n306);
   U51 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => O(9));
   U52 : AOI22_X1 port map( A1 => A0(9), A2 => n144, B1 => n178, B2 => A4(9), 
                           ZN => n310);
   U53 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161, 
                           C1 => A2(9), C2 => n153, ZN => n309);
   U54 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U55 : AOI22_X1 port map( A1 => A0(10), A2 => n139, B1 => A4(10), B2 => n178,
                           ZN => n185);
   U56 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => n156
                           , C1 => A2(10), C2 => n148, ZN => n184);
   U57 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U58 : AOI22_X1 port map( A1 => A0(11), A2 => n139, B1 => A4(11), B2 => n178,
                           ZN => n187);
   U59 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => n156
                           , C1 => A2(11), C2 => n148, ZN => n186);
   U60 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U61 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => n156
                           , C1 => A2(12), C2 => n148, ZN => n188);
   U62 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U63 : AOI22_X1 port map( A1 => A0(13), A2 => n139, B1 => A4(13), B2 => n177,
                           ZN => n191);
   U64 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => n156
                           , C1 => A2(13), C2 => n148, ZN => n190);
   U65 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U66 : AOI22_X1 port map( A1 => A0(14), A2 => n139, B1 => A4(14), B2 => n177,
                           ZN => n193);
   U67 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => n156
                           , C1 => A2(14), C2 => n148, ZN => n192);
   U68 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U69 : AOI22_X1 port map( A1 => A0(15), A2 => n139, B1 => A4(15), B2 => n177,
                           ZN => n195);
   U70 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n194);
   U71 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U72 : AOI22_X1 port map( A1 => A0(16), A2 => n139, B1 => A4(16), B2 => n177,
                           ZN => n197);
   U73 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n196);
   U74 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U75 : AOI22_X1 port map( A1 => A0(17), A2 => n139, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U76 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n198);
   U77 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U78 : AOI22_X1 port map( A1 => A0(18), A2 => n139, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U79 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => n156
                           , C1 => A2(18), C2 => n148, ZN => n200);
   U80 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U81 : AOI22_X1 port map( A1 => A0(25), A2 => n140, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U82 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => n157
                           , C1 => A2(25), C2 => n149, ZN => n216);
   U83 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U84 : AOI22_X1 port map( A1 => A0(19), A2 => n139, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U85 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n202);
   U86 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U87 : AOI22_X1 port map( A1 => A0(26), A2 => n140, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U88 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => n157
                           , C1 => A2(26), C2 => n149, ZN => n218);
   U89 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U90 : AOI22_X1 port map( A1 => A0(23), A2 => n140, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U91 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => n157
                           , C1 => A2(23), C2 => n149, ZN => n212);
   U92 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U93 : AOI22_X1 port map( A1 => A0(27), A2 => n140, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U94 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => n157
                           , C1 => A2(27), C2 => n149, ZN => n220);
   U95 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U96 : AOI22_X1 port map( A1 => A0(20), A2 => n140, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U97 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => n157
                           , C1 => A2(20), C2 => n149, ZN => n206);
   U98 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U99 : AOI22_X1 port map( A1 => A0(28), A2 => n140, B1 => A4(28), B2 => n176,
                           ZN => n223);
   U100 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => 
                           n157, C1 => A2(28), C2 => n149, ZN => n222);
   U101 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U102 : AOI22_X1 port map( A1 => A0(21), A2 => n140, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U103 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => 
                           n157, C1 => A2(21), C2 => n149, ZN => n208);
   U104 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U105 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => 
                           n157, C1 => A2(24), C2 => n149, ZN => n214);
   U106 : AOI22_X1 port map( A1 => A0(24), A2 => n140, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U107 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U108 : AOI22_X1 port map( A1 => A0(29), A2 => n140, B1 => A4(29), B2 => n176
                           , ZN => n225);
   U109 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => 
                           n157, C1 => A2(29), C2 => n149, ZN => n224);
   U110 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U111 : AOI22_X1 port map( A1 => A0(22), A2 => n140, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U112 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => 
                           n157, C1 => A2(22), C2 => n149, ZN => n210);
   U113 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U114 : AOI22_X1 port map( A1 => A0(30), A2 => n140, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U115 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => 
                           n157, C1 => A2(30), C2 => n149, ZN => n228);
   U116 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U117 : AOI22_X1 port map( A1 => A0(40), A2 => n141, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U118 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n250);
   U119 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U120 : AOI22_X1 port map( A1 => A0(31), A2 => n141, B1 => A4(31), B2 => n176
                           , ZN => n231);
   U121 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => 
                           n158, C1 => A2(31), C2 => n150, ZN => n230);
   U122 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U123 : AOI22_X1 port map( A1 => A0(32), A2 => n141, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U124 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => 
                           n158, C1 => A2(32), C2 => n150, ZN => n232);
   U125 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U126 : AOI22_X1 port map( A1 => A0(33), A2 => n141, B1 => A4(33), B2 => n176
                           , ZN => n235);
   U127 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => 
                           n158, C1 => A2(33), C2 => n150, ZN => n234);
   U128 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U129 : AOI22_X1 port map( A1 => A0(41), A2 => n141, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U130 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n252);
   U131 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U132 : AOI22_X1 port map( A1 => A0(34), A2 => n141, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U133 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n236);
   U134 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U135 : AOI22_X1 port map( A1 => A0(35), A2 => n141, B1 => A4(35), B2 => n175
                           , ZN => n239);
   U136 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n238);
   U137 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U138 : AOI22_X1 port map( A1 => A0(42), A2 => n142, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U139 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n254);
   U140 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U141 : AOI22_X1 port map( A1 => A0(36), A2 => n141, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U142 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n240);
   U143 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U144 : AOI22_X1 port map( A1 => A0(37), A2 => n141, B1 => A4(37), B2 => n175
                           , ZN => n243);
   U145 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n242);
   U146 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U147 : AOI22_X1 port map( A1 => A0(43), A2 => n142, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U148 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n256);
   U149 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U150 : AOI22_X1 port map( A1 => A0(38), A2 => n141, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U151 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n244);
   U152 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U153 : AOI22_X1 port map( A1 => A0(39), A2 => n141, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U154 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => 
                           n158, C1 => A2(39), C2 => n150, ZN => n246);
   U155 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U156 : AOI22_X1 port map( A1 => A0(44), A2 => n142, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U157 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n258);
   U158 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U159 : AOI22_X1 port map( A1 => A0(45), A2 => n142, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U160 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n260);
   U161 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U162 : AOI22_X1 port map( A1 => A0(46), A2 => n142, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U163 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n262);
   U164 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U165 : AOI22_X1 port map( A1 => A0(47), A2 => n142, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U166 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n264);
   U167 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U168 : AOI22_X1 port map( A1 => A0(48), A2 => n142, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U169 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n266);
   U170 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U171 : AOI22_X1 port map( A1 => A0(49), A2 => n142, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U172 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n268);
   U173 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U174 : AOI22_X1 port map( A1 => A0(50), A2 => n142, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U175 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n272);
   U176 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U177 : AOI22_X1 port map( A1 => A0(51), A2 => n142, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U178 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n274);
   U179 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U180 : AOI22_X1 port map( A1 => A0(52), A2 => n142, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U181 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n276);
   U182 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U183 : AOI22_X1 port map( A1 => A0(53), A2 => n143, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U184 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n278);
   U185 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U186 : AOI22_X1 port map( A1 => A0(54), A2 => n143, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U187 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n280);
   U188 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U189 : AOI22_X1 port map( A1 => A0(55), A2 => n143, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U190 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n282);
   U191 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U192 : AOI22_X1 port map( A1 => A0(56), A2 => n143, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U193 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n284);
   U194 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U195 : AOI22_X1 port map( A1 => A0(57), A2 => n143, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U196 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n286);
   U197 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U198 : AOI22_X1 port map( A1 => A0(58), A2 => n143, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U199 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n288);
   U200 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U201 : AOI22_X1 port map( A1 => A0(59), A2 => n143, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U202 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n290);
   U203 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U204 : AOI22_X1 port map( A1 => A0(60), A2 => n143, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U205 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n294);
   U206 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U207 : AOI22_X1 port map( A1 => A0(61), A2 => n143, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U208 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n296);
   U209 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U210 : AOI22_X1 port map( A1 => A0(62), A2 => n143, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U211 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n298);
   U212 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U213 : AOI22_X1 port map( A1 => A0(63), A2 => n143, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U214 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n300);
   U215 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U216 : AOI22_X1 port map( A1 => A0(0), A2 => n139, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U217 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n182);
   U218 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U219 : AOI22_X1 port map( A1 => A0(1), A2 => n139, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U220 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n204);
   U221 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U222 : AOI22_X1 port map( A1 => A0(2), A2 => n140, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U223 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n226);
   U224 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U225 : AOI22_X1 port map( A1 => A0(3), A2 => n141, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U226 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n248);
   U227 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U228 : AOI22_X1 port map( A1 => A0(4), A2 => n142, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U229 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n270);
   U230 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U231 : AOI22_X1 port map( A1 => A0(5), A2 => n143, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U232 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n292);
   U233 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U234 : AOI22_X1 port map( A1 => A0(6), A2 => n144, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U235 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161,
                           C1 => A2(6), C2 => n153, ZN => n302);
   U236 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U237 : AOI22_X1 port map( A1 => A0(7), A2 => n144, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U238 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161,
                           C1 => A2(7), C2 => n153, ZN => n304);
   U239 : AOI22_X1 port map( A1 => A0(12), A2 => n139, B1 => A4(12), B2 => n177
                           , ZN => n189);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_11 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_11;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n136, Z => n154);
   U2 : CLKBUF_X1 port map( A => n138, Z => n162);
   U3 : CLKBUF_X1 port map( A => n137, Z => n170);
   U4 : CLKBUF_X1 port map( A => n172, Z => n180);
   U5 : BUF_X1 port map( A => n136, Z => n155);
   U6 : BUF_X1 port map( A => n137, Z => n171);
   U7 : BUF_X1 port map( A => n138, Z => n163);
   U8 : BUF_X1 port map( A => n147, Z => n146);
   U9 : BUF_X1 port map( A => n147, Z => n145);
   U10 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U11 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n137);
   U12 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U13 : BUF_X1 port map( A => n172, Z => n179);
   U14 : BUF_X1 port map( A => sel(2), Z => n172);
   U15 : BUF_X1 port map( A => n155, Z => n148);
   U16 : BUF_X1 port map( A => n171, Z => n164);
   U17 : BUF_X1 port map( A => n163, Z => n156);
   U18 : BUF_X1 port map( A => n171, Z => n165);
   U19 : BUF_X1 port map( A => n155, Z => n149);
   U20 : BUF_X1 port map( A => n163, Z => n157);
   U21 : BUF_X1 port map( A => n171, Z => n166);
   U22 : BUF_X1 port map( A => n155, Z => n150);
   U23 : BUF_X1 port map( A => n163, Z => n158);
   U24 : BUF_X1 port map( A => n170, Z => n167);
   U25 : BUF_X1 port map( A => n154, Z => n151);
   U26 : BUF_X1 port map( A => n162, Z => n159);
   U27 : BUF_X1 port map( A => n170, Z => n168);
   U28 : BUF_X1 port map( A => n154, Z => n152);
   U29 : BUF_X1 port map( A => n162, Z => n160);
   U30 : BUF_X1 port map( A => n146, Z => n140);
   U31 : BUF_X1 port map( A => n146, Z => n141);
   U32 : BUF_X1 port map( A => n145, Z => n142);
   U33 : BUF_X1 port map( A => n145, Z => n143);
   U34 : BUF_X1 port map( A => n146, Z => n139);
   U35 : BUF_X1 port map( A => n145, Z => n144);
   U36 : BUF_X1 port map( A => n162, Z => n161);
   U37 : BUF_X1 port map( A => n154, Z => n153);
   U38 : BUF_X1 port map( A => n170, Z => n169);
   U39 : BUF_X1 port map( A => n179, Z => n178);
   U40 : BUF_X1 port map( A => n179, Z => n177);
   U41 : BUF_X1 port map( A => n179, Z => n176);
   U42 : BUF_X1 port map( A => n180, Z => n175);
   U43 : BUF_X1 port map( A => n180, Z => n174);
   U44 : BUF_X1 port map( A => n180, Z => n173);
   U45 : INV_X1 port map( A => sel(0), ZN => n181);
   U46 : BUF_X1 port map( A => n308, Z => n147);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U49 : AOI22_X1 port map( A1 => A0(10), A2 => n139, B1 => A4(10), B2 => n178,
                           ZN => n185);
   U50 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => n156
                           , C1 => A2(10), C2 => n148, ZN => n184);
   U51 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U52 : AOI22_X1 port map( A1 => A0(11), A2 => n139, B1 => A4(11), B2 => n178,
                           ZN => n187);
   U53 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => n156
                           , C1 => A2(11), C2 => n148, ZN => n186);
   U54 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U55 : AOI22_X1 port map( A1 => A0(12), A2 => n139, B1 => A4(12), B2 => n177,
                           ZN => n189);
   U56 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => n156
                           , C1 => A2(12), C2 => n148, ZN => n188);
   U57 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U58 : AOI22_X1 port map( A1 => A0(13), A2 => n139, B1 => A4(13), B2 => n177,
                           ZN => n191);
   U59 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => n156
                           , C1 => A2(13), C2 => n148, ZN => n190);
   U60 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U61 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => n156
                           , C1 => A2(14), C2 => n148, ZN => n192);
   U62 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U63 : AOI22_X1 port map( A1 => A0(15), A2 => n139, B1 => A4(15), B2 => n177,
                           ZN => n195);
   U64 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n194);
   U65 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U66 : AOI22_X1 port map( A1 => A0(16), A2 => n139, B1 => A4(16), B2 => n177,
                           ZN => n197);
   U67 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n196);
   U68 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U69 : AOI22_X1 port map( A1 => A0(17), A2 => n139, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U70 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n198);
   U71 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U72 : AOI22_X1 port map( A1 => A0(18), A2 => n139, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U73 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => n156
                           , C1 => A2(18), C2 => n148, ZN => n200);
   U74 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U75 : AOI22_X1 port map( A1 => A0(19), A2 => n139, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U76 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n202);
   U77 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U78 : AOI22_X1 port map( A1 => A0(20), A2 => n140, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U79 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => n157
                           , C1 => A2(20), C2 => n149, ZN => n206);
   U80 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U81 : AOI22_X1 port map( A1 => A0(27), A2 => n140, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U82 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => n157
                           , C1 => A2(27), C2 => n149, ZN => n220);
   U83 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U84 : AOI22_X1 port map( A1 => A0(21), A2 => n140, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U85 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => n157
                           , C1 => A2(21), C2 => n149, ZN => n208);
   U86 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U87 : AOI22_X1 port map( A1 => A0(28), A2 => n140, B1 => A4(28), B2 => n176,
                           ZN => n223);
   U88 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => n157
                           , C1 => A2(28), C2 => n149, ZN => n222);
   U89 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U90 : AOI22_X1 port map( A1 => A0(25), A2 => n140, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U91 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => n157
                           , C1 => A2(25), C2 => n149, ZN => n216);
   U92 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U93 : AOI22_X1 port map( A1 => A0(29), A2 => n140, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U94 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => n157
                           , C1 => A2(29), C2 => n149, ZN => n224);
   U95 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U96 : AOI22_X1 port map( A1 => A0(22), A2 => n140, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U97 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => n157
                           , C1 => A2(22), C2 => n149, ZN => n210);
   U98 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U99 : AOI22_X1 port map( A1 => A0(30), A2 => n140, B1 => A4(30), B2 => n176,
                           ZN => n229);
   U100 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => 
                           n157, C1 => A2(30), C2 => n149, ZN => n228);
   U101 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U102 : AOI22_X1 port map( A1 => A0(23), A2 => n140, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U103 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => 
                           n157, C1 => A2(23), C2 => n149, ZN => n212);
   U104 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U105 : AOI22_X1 port map( A1 => A0(31), A2 => n141, B1 => A4(31), B2 => n176
                           , ZN => n231);
   U106 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => 
                           n158, C1 => A2(31), C2 => n150, ZN => n230);
   U107 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U108 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => 
                           n157, C1 => A2(26), C2 => n149, ZN => n218);
   U109 : AOI22_X1 port map( A1 => A0(26), A2 => n140, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U110 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U111 : AOI22_X1 port map( A1 => A0(24), A2 => n140, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U112 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => 
                           n157, C1 => A2(24), C2 => n149, ZN => n214);
   U113 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U114 : AOI22_X1 port map( A1 => A0(32), A2 => n141, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U115 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => 
                           n158, C1 => A2(32), C2 => n150, ZN => n232);
   U116 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U117 : AOI22_X1 port map( A1 => A0(33), A2 => n141, B1 => A4(33), B2 => n176
                           , ZN => n235);
   U118 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => 
                           n158, C1 => A2(33), C2 => n150, ZN => n234);
   U119 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U120 : AOI22_X1 port map( A1 => A0(42), A2 => n142, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U121 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n254);
   U122 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U123 : AOI22_X1 port map( A1 => A0(34), A2 => n141, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U124 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n236);
   U125 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U126 : AOI22_X1 port map( A1 => A0(35), A2 => n141, B1 => A4(35), B2 => n175
                           , ZN => n239);
   U127 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n238);
   U128 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U129 : AOI22_X1 port map( A1 => A0(43), A2 => n142, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U130 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n256);
   U131 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U132 : AOI22_X1 port map( A1 => A0(36), A2 => n141, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U133 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n240);
   U134 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U135 : AOI22_X1 port map( A1 => A0(37), A2 => n141, B1 => A4(37), B2 => n175
                           , ZN => n243);
   U136 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n242);
   U137 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U138 : AOI22_X1 port map( A1 => A0(44), A2 => n142, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U139 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n258);
   U140 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U141 : AOI22_X1 port map( A1 => A0(38), A2 => n141, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U142 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n244);
   U143 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U144 : AOI22_X1 port map( A1 => A0(39), A2 => n141, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U145 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => 
                           n158, C1 => A2(39), C2 => n150, ZN => n246);
   U146 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U147 : AOI22_X1 port map( A1 => A0(40), A2 => n141, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U148 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n250);
   U149 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U150 : AOI22_X1 port map( A1 => A0(45), A2 => n142, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U151 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n260);
   U152 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U153 : AOI22_X1 port map( A1 => A0(41), A2 => n141, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U154 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n252);
   U155 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U156 : AOI22_X1 port map( A1 => A0(46), A2 => n142, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U157 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n262);
   U158 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U159 : AOI22_X1 port map( A1 => A0(47), A2 => n142, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U160 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n264);
   U161 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U162 : AOI22_X1 port map( A1 => A0(48), A2 => n142, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U163 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n266);
   U164 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U165 : AOI22_X1 port map( A1 => A0(49), A2 => n142, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U166 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n268);
   U167 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U168 : AOI22_X1 port map( A1 => A0(50), A2 => n142, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U169 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n272);
   U170 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U171 : AOI22_X1 port map( A1 => A0(51), A2 => n142, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U172 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n274);
   U173 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U174 : AOI22_X1 port map( A1 => A0(52), A2 => n142, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U175 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n276);
   U176 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U177 : AOI22_X1 port map( A1 => A0(53), A2 => n143, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U178 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n278);
   U179 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U180 : AOI22_X1 port map( A1 => A0(54), A2 => n143, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U181 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n280);
   U182 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U183 : AOI22_X1 port map( A1 => A0(55), A2 => n143, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U184 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n282);
   U185 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U186 : AOI22_X1 port map( A1 => A0(56), A2 => n143, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U187 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n284);
   U188 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U189 : AOI22_X1 port map( A1 => A0(57), A2 => n143, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U190 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n286);
   U191 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U192 : AOI22_X1 port map( A1 => A0(58), A2 => n143, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U193 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n288);
   U194 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U195 : AOI22_X1 port map( A1 => A0(59), A2 => n143, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U196 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n290);
   U197 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U198 : AOI22_X1 port map( A1 => A0(60), A2 => n143, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U199 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n294);
   U200 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U201 : AOI22_X1 port map( A1 => A0(61), A2 => n143, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U202 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n296);
   U203 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U204 : AOI22_X1 port map( A1 => A0(62), A2 => n143, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U205 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n298);
   U206 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U207 : AOI22_X1 port map( A1 => A0(63), A2 => n143, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U208 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n300);
   U209 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U210 : AOI22_X1 port map( A1 => A0(0), A2 => n139, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U211 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n182);
   U212 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U213 : AOI22_X1 port map( A1 => A0(1), A2 => n139, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U214 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n204);
   U215 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U216 : AOI22_X1 port map( A1 => A0(2), A2 => n140, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U217 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n226);
   U218 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U219 : AOI22_X1 port map( A1 => A0(3), A2 => n141, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U220 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n248);
   U221 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U222 : AOI22_X1 port map( A1 => A0(4), A2 => n142, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U223 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n270);
   U224 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U225 : AOI22_X1 port map( A1 => A0(5), A2 => n143, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U226 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n292);
   U227 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U228 : AOI22_X1 port map( A1 => A0(6), A2 => n144, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U229 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161,
                           C1 => A2(6), C2 => n153, ZN => n302);
   U230 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U231 : AOI22_X1 port map( A1 => A0(7), A2 => n144, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U232 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161,
                           C1 => A2(7), C2 => n153, ZN => n304);
   U233 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U234 : AOI22_X1 port map( A1 => A0(8), A2 => n144, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U235 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161,
                           C1 => A2(8), C2 => n153, ZN => n306);
   U236 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => O(9));
   U237 : AOI22_X1 port map( A1 => A0(9), A2 => n144, B1 => n178, B2 => A4(9), 
                           ZN => n310);
   U238 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161,
                           C1 => A2(9), C2 => n153, ZN => n309);
   U239 : AOI22_X1 port map( A1 => A0(14), A2 => n139, B1 => A4(14), B2 => n177
                           , ZN => n193);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_10 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_10;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n136, Z => n155);
   U2 : BUF_X1 port map( A => n137, Z => n171);
   U3 : BUF_X1 port map( A => n138, Z => n163);
   U4 : BUF_X1 port map( A => n136, Z => n154);
   U5 : BUF_X1 port map( A => n137, Z => n170);
   U6 : BUF_X1 port map( A => n138, Z => n162);
   U7 : BUF_X1 port map( A => n147, Z => n146);
   U8 : BUF_X1 port map( A => n147, Z => n145);
   U9 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U10 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n137);
   U11 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U12 : BUF_X1 port map( A => n172, Z => n179);
   U13 : BUF_X1 port map( A => n172, Z => n180);
   U14 : BUF_X1 port map( A => sel(2), Z => n172);
   U15 : BUF_X1 port map( A => n155, Z => n148);
   U16 : BUF_X1 port map( A => n171, Z => n164);
   U17 : BUF_X1 port map( A => n163, Z => n156);
   U18 : BUF_X1 port map( A => n171, Z => n165);
   U19 : BUF_X1 port map( A => n155, Z => n149);
   U20 : BUF_X1 port map( A => n163, Z => n157);
   U21 : BUF_X1 port map( A => n171, Z => n166);
   U22 : BUF_X1 port map( A => n155, Z => n150);
   U23 : BUF_X1 port map( A => n163, Z => n158);
   U24 : BUF_X1 port map( A => n170, Z => n167);
   U25 : BUF_X1 port map( A => n154, Z => n151);
   U26 : BUF_X1 port map( A => n162, Z => n159);
   U27 : BUF_X1 port map( A => n170, Z => n168);
   U28 : BUF_X1 port map( A => n154, Z => n152);
   U29 : BUF_X1 port map( A => n162, Z => n160);
   U30 : BUF_X1 port map( A => n146, Z => n140);
   U31 : BUF_X1 port map( A => n146, Z => n141);
   U32 : BUF_X1 port map( A => n145, Z => n142);
   U33 : BUF_X1 port map( A => n145, Z => n143);
   U34 : BUF_X1 port map( A => n146, Z => n139);
   U35 : BUF_X1 port map( A => n145, Z => n144);
   U36 : BUF_X1 port map( A => n162, Z => n161);
   U37 : BUF_X1 port map( A => n154, Z => n153);
   U38 : BUF_X1 port map( A => n170, Z => n169);
   U39 : BUF_X1 port map( A => n179, Z => n177);
   U40 : BUF_X1 port map( A => n179, Z => n176);
   U41 : BUF_X1 port map( A => n180, Z => n175);
   U42 : BUF_X1 port map( A => n180, Z => n174);
   U43 : BUF_X1 port map( A => n180, Z => n173);
   U44 : BUF_X1 port map( A => n179, Z => n178);
   U45 : INV_X1 port map( A => sel(0), ZN => n181);
   U46 : BUF_X1 port map( A => n308, Z => n147);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U49 : AOI22_X1 port map( A1 => A0(12), A2 => n139, B1 => A4(12), B2 => n177,
                           ZN => n189);
   U50 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => n156
                           , C1 => A2(12), C2 => n148, ZN => n188);
   U51 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U52 : AOI22_X1 port map( A1 => A0(13), A2 => n139, B1 => A4(13), B2 => n177,
                           ZN => n191);
   U53 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => n156
                           , C1 => A2(13), C2 => n148, ZN => n190);
   U54 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U55 : AOI22_X1 port map( A1 => A0(14), A2 => n139, B1 => A4(14), B2 => n177,
                           ZN => n193);
   U56 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => n156
                           , C1 => A2(14), C2 => n148, ZN => n192);
   U57 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U58 : AOI22_X1 port map( A1 => A0(15), A2 => n139, B1 => A4(15), B2 => n177,
                           ZN => n195);
   U59 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n194);
   U60 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U61 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n196);
   U62 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U63 : AOI22_X1 port map( A1 => A0(17), A2 => n139, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U64 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n198);
   U65 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U66 : AOI22_X1 port map( A1 => A0(18), A2 => n139, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U67 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => n156
                           , C1 => A2(18), C2 => n148, ZN => n200);
   U68 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U69 : AOI22_X1 port map( A1 => A0(19), A2 => n139, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U70 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n202);
   U71 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U72 : AOI22_X1 port map( A1 => A0(20), A2 => n140, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U73 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => n157
                           , C1 => A2(20), C2 => n149, ZN => n206);
   U74 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U75 : AOI22_X1 port map( A1 => A0(21), A2 => n140, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U76 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => n157
                           , C1 => A2(21), C2 => n149, ZN => n208);
   U77 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U78 : AOI22_X1 port map( A1 => A0(22), A2 => n140, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U79 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => n157
                           , C1 => A2(22), C2 => n149, ZN => n210);
   U80 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U81 : AOI22_X1 port map( A1 => A0(29), A2 => n140, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U82 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => n157
                           , C1 => A2(29), C2 => n149, ZN => n224);
   U83 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U84 : AOI22_X1 port map( A1 => A0(30), A2 => n140, B1 => A4(30), B2 => n176,
                           ZN => n229);
   U85 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => n157
                           , C1 => A2(30), C2 => n149, ZN => n228);
   U86 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U87 : AOI22_X1 port map( A1 => A0(27), A2 => n140, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U88 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => n157
                           , C1 => A2(27), C2 => n149, ZN => n220);
   U89 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U90 : AOI22_X1 port map( A1 => A0(23), A2 => n140, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U91 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => n157
                           , C1 => A2(23), C2 => n149, ZN => n212);
   U92 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U93 : AOI22_X1 port map( A1 => A0(31), A2 => n141, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U94 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => n158
                           , C1 => A2(31), C2 => n150, ZN => n230);
   U95 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U96 : AOI22_X1 port map( A1 => A0(24), A2 => n140, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U97 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => n157
                           , C1 => A2(24), C2 => n149, ZN => n214);
   U98 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U99 : AOI22_X1 port map( A1 => A0(32), A2 => n141, B1 => A4(32), B2 => n176,
                           ZN => n233);
   U100 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => 
                           n158, C1 => A2(32), C2 => n150, ZN => n232);
   U101 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U102 : AOI22_X1 port map( A1 => A0(25), A2 => n140, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U103 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => 
                           n157, C1 => A2(25), C2 => n149, ZN => n216);
   U104 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U105 : AOI22_X1 port map( A1 => A0(33), A2 => n141, B1 => A4(33), B2 => n176
                           , ZN => n235);
   U106 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => 
                           n158, C1 => A2(33), C2 => n150, ZN => n234);
   U107 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U108 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => 
                           n157, C1 => A2(28), C2 => n149, ZN => n222);
   U109 : AOI22_X1 port map( A1 => A0(28), A2 => n140, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U110 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U111 : AOI22_X1 port map( A1 => A0(26), A2 => n140, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U112 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => 
                           n157, C1 => A2(26), C2 => n149, ZN => n218);
   U113 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U114 : AOI22_X1 port map( A1 => A0(34), A2 => n141, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U115 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n236);
   U116 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U117 : AOI22_X1 port map( A1 => A0(35), A2 => n141, B1 => A4(35), B2 => n175
                           , ZN => n239);
   U118 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n238);
   U119 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U120 : AOI22_X1 port map( A1 => A0(44), A2 => n142, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U121 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n258);
   U122 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U123 : AOI22_X1 port map( A1 => A0(36), A2 => n141, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U124 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n240);
   U125 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U126 : AOI22_X1 port map( A1 => A0(37), A2 => n141, B1 => A4(37), B2 => n175
                           , ZN => n243);
   U127 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n242);
   U128 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U129 : AOI22_X1 port map( A1 => A0(45), A2 => n142, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U130 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n260);
   U131 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U132 : AOI22_X1 port map( A1 => A0(38), A2 => n141, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U133 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n244);
   U134 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U135 : AOI22_X1 port map( A1 => A0(39), A2 => n141, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U136 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => 
                           n158, C1 => A2(39), C2 => n150, ZN => n246);
   U137 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U138 : AOI22_X1 port map( A1 => A0(46), A2 => n142, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U139 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n262);
   U140 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U141 : AOI22_X1 port map( A1 => A0(40), A2 => n141, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U142 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n250);
   U143 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U144 : AOI22_X1 port map( A1 => A0(41), A2 => n141, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U145 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n252);
   U146 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U147 : AOI22_X1 port map( A1 => A0(47), A2 => n142, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U148 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n264);
   U149 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U150 : AOI22_X1 port map( A1 => A0(42), A2 => n142, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U151 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n254);
   U152 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U153 : AOI22_X1 port map( A1 => A0(43), A2 => n142, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U154 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n256);
   U155 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U156 : AOI22_X1 port map( A1 => A0(48), A2 => n142, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U157 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n266);
   U158 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U159 : AOI22_X1 port map( A1 => A0(49), A2 => n142, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U160 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n268);
   U161 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U162 : AOI22_X1 port map( A1 => A0(50), A2 => n142, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U163 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n272);
   U164 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U165 : AOI22_X1 port map( A1 => A0(51), A2 => n142, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U166 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n274);
   U167 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U168 : AOI22_X1 port map( A1 => A0(52), A2 => n142, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U169 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n276);
   U170 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U171 : AOI22_X1 port map( A1 => A0(53), A2 => n143, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U172 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n278);
   U173 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U174 : AOI22_X1 port map( A1 => A0(54), A2 => n143, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U175 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n280);
   U176 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U177 : AOI22_X1 port map( A1 => A0(55), A2 => n143, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U178 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n282);
   U179 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U180 : AOI22_X1 port map( A1 => A0(56), A2 => n143, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U181 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n284);
   U182 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U183 : AOI22_X1 port map( A1 => A0(57), A2 => n143, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U184 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n286);
   U185 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U186 : AOI22_X1 port map( A1 => A0(58), A2 => n143, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U187 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n288);
   U188 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U189 : AOI22_X1 port map( A1 => A0(59), A2 => n143, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U190 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n290);
   U191 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U192 : AOI22_X1 port map( A1 => A0(60), A2 => n143, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U193 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n294);
   U194 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U195 : AOI22_X1 port map( A1 => A0(61), A2 => n143, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U196 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n296);
   U197 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U198 : AOI22_X1 port map( A1 => A0(62), A2 => n143, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U199 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n298);
   U200 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U201 : AOI22_X1 port map( A1 => A0(63), A2 => n143, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U202 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n300);
   U203 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U204 : AOI22_X1 port map( A1 => A0(0), A2 => n139, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U205 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n182);
   U206 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U207 : AOI22_X1 port map( A1 => A0(1), A2 => n139, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U208 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n204);
   U209 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U210 : AOI22_X1 port map( A1 => A0(2), A2 => n140, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U211 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n226);
   U212 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U213 : AOI22_X1 port map( A1 => A0(3), A2 => n141, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U214 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n248);
   U215 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U216 : AOI22_X1 port map( A1 => A0(4), A2 => n142, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U217 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n270);
   U218 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U219 : AOI22_X1 port map( A1 => A0(5), A2 => n143, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U220 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n292);
   U221 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U222 : AOI22_X1 port map( A1 => A0(6), A2 => n144, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U223 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161,
                           C1 => A2(6), C2 => n153, ZN => n302);
   U224 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U225 : AOI22_X1 port map( A1 => A0(7), A2 => n144, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U226 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161,
                           C1 => A2(7), C2 => n153, ZN => n304);
   U227 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U228 : AOI22_X1 port map( A1 => A0(8), A2 => n144, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U229 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161,
                           C1 => A2(8), C2 => n153, ZN => n306);
   U230 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => O(9));
   U231 : AOI22_X1 port map( A1 => A0(9), A2 => n144, B1 => n178, B2 => A4(9), 
                           ZN => n310);
   U232 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161,
                           C1 => A2(9), C2 => n153, ZN => n309);
   U233 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U234 : AOI22_X1 port map( A1 => A0(10), A2 => n139, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U235 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => 
                           n156, C1 => A2(10), C2 => n148, ZN => n184);
   U236 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U237 : AOI22_X1 port map( A1 => A0(11), A2 => n139, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U238 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => 
                           n156, C1 => A2(11), C2 => n148, ZN => n186);
   U239 : AOI22_X1 port map( A1 => A0(16), A2 => n139, B1 => A4(16), B2 => n177
                           , ZN => n197);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_9 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_9;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n136, Z => n155);
   U2 : BUF_X1 port map( A => n137, Z => n171);
   U3 : BUF_X1 port map( A => n138, Z => n163);
   U4 : BUF_X1 port map( A => n136, Z => n154);
   U5 : BUF_X1 port map( A => n137, Z => n170);
   U6 : BUF_X1 port map( A => n138, Z => n162);
   U7 : BUF_X1 port map( A => n147, Z => n146);
   U8 : BUF_X1 port map( A => n147, Z => n145);
   U9 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U10 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n137);
   U11 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n138);
   U12 : BUF_X1 port map( A => n172, Z => n179);
   U13 : BUF_X1 port map( A => n172, Z => n180);
   U14 : BUF_X1 port map( A => sel(2), Z => n172);
   U15 : BUF_X1 port map( A => n155, Z => n148);
   U16 : BUF_X1 port map( A => n171, Z => n164);
   U17 : BUF_X1 port map( A => n163, Z => n156);
   U18 : BUF_X1 port map( A => n171, Z => n165);
   U19 : BUF_X1 port map( A => n155, Z => n149);
   U20 : BUF_X1 port map( A => n163, Z => n157);
   U21 : BUF_X1 port map( A => n171, Z => n166);
   U22 : BUF_X1 port map( A => n155, Z => n150);
   U23 : BUF_X1 port map( A => n163, Z => n158);
   U24 : BUF_X1 port map( A => n170, Z => n167);
   U25 : BUF_X1 port map( A => n154, Z => n151);
   U26 : BUF_X1 port map( A => n162, Z => n159);
   U27 : BUF_X1 port map( A => n170, Z => n168);
   U28 : BUF_X1 port map( A => n154, Z => n152);
   U29 : BUF_X1 port map( A => n162, Z => n160);
   U30 : BUF_X1 port map( A => n146, Z => n140);
   U31 : BUF_X1 port map( A => n146, Z => n141);
   U32 : BUF_X1 port map( A => n145, Z => n142);
   U33 : BUF_X1 port map( A => n145, Z => n143);
   U34 : BUF_X1 port map( A => n146, Z => n139);
   U35 : BUF_X1 port map( A => n145, Z => n144);
   U36 : BUF_X1 port map( A => n162, Z => n161);
   U37 : BUF_X1 port map( A => n154, Z => n153);
   U38 : BUF_X1 port map( A => n170, Z => n169);
   U39 : BUF_X1 port map( A => n179, Z => n177);
   U40 : BUF_X1 port map( A => n179, Z => n176);
   U41 : BUF_X1 port map( A => n180, Z => n175);
   U42 : BUF_X1 port map( A => n180, Z => n174);
   U43 : BUF_X1 port map( A => n180, Z => n173);
   U44 : BUF_X1 port map( A => n179, Z => n178);
   U45 : INV_X1 port map( A => sel(0), ZN => n181);
   U46 : BUF_X1 port map( A => n308, Z => n147);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U49 : AOI22_X1 port map( A1 => A0(14), A2 => n139, B1 => A4(14), B2 => n177,
                           ZN => n193);
   U50 : AOI222_X1 port map( A1 => A1(14), A2 => n164, B1 => A3(14), B2 => n156
                           , C1 => A2(14), C2 => n148, ZN => n192);
   U51 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U52 : AOI22_X1 port map( A1 => A0(15), A2 => n139, B1 => A4(15), B2 => n177,
                           ZN => n195);
   U53 : AOI222_X1 port map( A1 => A1(15), A2 => n164, B1 => A3(15), B2 => n156
                           , C1 => A2(15), C2 => n148, ZN => n194);
   U54 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U55 : AOI22_X1 port map( A1 => A0(16), A2 => n139, B1 => A4(16), B2 => n177,
                           ZN => n197);
   U56 : AOI222_X1 port map( A1 => A1(16), A2 => n164, B1 => A3(16), B2 => n156
                           , C1 => A2(16), C2 => n148, ZN => n196);
   U57 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U58 : AOI22_X1 port map( A1 => A0(17), A2 => n139, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U59 : AOI222_X1 port map( A1 => A1(17), A2 => n164, B1 => A3(17), B2 => n156
                           , C1 => A2(17), C2 => n148, ZN => n198);
   U60 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U61 : AOI222_X1 port map( A1 => A1(18), A2 => n164, B1 => A3(18), B2 => n156
                           , C1 => A2(18), C2 => n148, ZN => n200);
   U62 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U63 : AOI22_X1 port map( A1 => A0(19), A2 => n139, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U64 : AOI222_X1 port map( A1 => A1(19), A2 => n164, B1 => A3(19), B2 => n156
                           , C1 => A2(19), C2 => n148, ZN => n202);
   U65 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U66 : AOI22_X1 port map( A1 => A0(20), A2 => n140, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U67 : AOI222_X1 port map( A1 => A1(20), A2 => n165, B1 => A3(20), B2 => n157
                           , C1 => A2(20), C2 => n149, ZN => n206);
   U68 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U69 : AOI22_X1 port map( A1 => A0(21), A2 => n140, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U70 : AOI222_X1 port map( A1 => A1(21), A2 => n165, B1 => A3(21), B2 => n157
                           , C1 => A2(21), C2 => n149, ZN => n208);
   U71 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U72 : AOI22_X1 port map( A1 => A0(22), A2 => n140, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U73 : AOI222_X1 port map( A1 => A1(22), A2 => n165, B1 => A3(22), B2 => n157
                           , C1 => A2(22), C2 => n149, ZN => n210);
   U74 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U75 : AOI22_X1 port map( A1 => A0(23), A2 => n140, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U76 : AOI222_X1 port map( A1 => A1(23), A2 => n165, B1 => A3(23), B2 => n157
                           , C1 => A2(23), C2 => n149, ZN => n212);
   U77 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U78 : AOI22_X1 port map( A1 => A0(24), A2 => n140, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U79 : AOI222_X1 port map( A1 => A1(24), A2 => n165, B1 => A3(24), B2 => n157
                           , C1 => A2(24), C2 => n149, ZN => n214);
   U80 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U81 : AOI22_X1 port map( A1 => A0(31), A2 => n141, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U82 : AOI222_X1 port map( A1 => A1(31), A2 => n166, B1 => A3(31), B2 => n158
                           , C1 => A2(31), C2 => n150, ZN => n230);
   U83 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U84 : AOI22_X1 port map( A1 => A0(32), A2 => n141, B1 => A4(32), B2 => n176,
                           ZN => n233);
   U85 : AOI222_X1 port map( A1 => A1(32), A2 => n166, B1 => A3(32), B2 => n158
                           , C1 => A2(32), C2 => n150, ZN => n232);
   U86 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U87 : AOI22_X1 port map( A1 => A0(29), A2 => n140, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U88 : AOI222_X1 port map( A1 => A1(29), A2 => n165, B1 => A3(29), B2 => n157
                           , C1 => A2(29), C2 => n149, ZN => n224);
   U89 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U90 : AOI22_X1 port map( A1 => A0(25), A2 => n140, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U91 : AOI222_X1 port map( A1 => A1(25), A2 => n165, B1 => A3(25), B2 => n157
                           , C1 => A2(25), C2 => n149, ZN => n216);
   U92 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U93 : AOI22_X1 port map( A1 => A0(33), A2 => n141, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U94 : AOI222_X1 port map( A1 => A1(33), A2 => n166, B1 => A3(33), B2 => n158
                           , C1 => A2(33), C2 => n150, ZN => n234);
   U95 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U96 : AOI22_X1 port map( A1 => A0(26), A2 => n140, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U97 : AOI222_X1 port map( A1 => A1(26), A2 => n165, B1 => A3(26), B2 => n157
                           , C1 => A2(26), C2 => n149, ZN => n218);
   U98 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U99 : AOI22_X1 port map( A1 => A0(34), A2 => n141, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U100 : AOI222_X1 port map( A1 => A1(34), A2 => n166, B1 => A3(34), B2 => 
                           n158, C1 => A2(34), C2 => n150, ZN => n236);
   U101 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U102 : AOI22_X1 port map( A1 => A0(27), A2 => n140, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U103 : AOI222_X1 port map( A1 => A1(27), A2 => n165, B1 => A3(27), B2 => 
                           n157, C1 => A2(27), C2 => n149, ZN => n220);
   U104 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U105 : AOI22_X1 port map( A1 => A0(35), A2 => n141, B1 => A4(35), B2 => n175
                           , ZN => n239);
   U106 : AOI222_X1 port map( A1 => A1(35), A2 => n166, B1 => A3(35), B2 => 
                           n158, C1 => A2(35), C2 => n150, ZN => n238);
   U107 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U108 : AOI22_X1 port map( A1 => A0(28), A2 => n140, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U109 : AOI222_X1 port map( A1 => A1(28), A2 => n165, B1 => A3(28), B2 => 
                           n157, C1 => A2(28), C2 => n149, ZN => n222);
   U110 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U111 : AOI222_X1 port map( A1 => A1(30), A2 => n165, B1 => A3(30), B2 => 
                           n157, C1 => A2(30), C2 => n149, ZN => n228);
   U112 : AOI22_X1 port map( A1 => A0(30), A2 => n140, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U113 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U114 : AOI22_X1 port map( A1 => A0(36), A2 => n141, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U115 : AOI222_X1 port map( A1 => A1(36), A2 => n166, B1 => A3(36), B2 => 
                           n158, C1 => A2(36), C2 => n150, ZN => n240);
   U116 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U117 : AOI22_X1 port map( A1 => A0(37), A2 => n141, B1 => A4(37), B2 => n175
                           , ZN => n243);
   U118 : AOI222_X1 port map( A1 => A1(37), A2 => n166, B1 => A3(37), B2 => 
                           n158, C1 => A2(37), C2 => n150, ZN => n242);
   U119 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U120 : AOI22_X1 port map( A1 => A0(46), A2 => n142, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U121 : AOI222_X1 port map( A1 => A1(46), A2 => n167, B1 => A3(46), B2 => 
                           n159, C1 => A2(46), C2 => n151, ZN => n262);
   U122 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U123 : AOI22_X1 port map( A1 => A0(38), A2 => n141, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U124 : AOI222_X1 port map( A1 => A1(38), A2 => n166, B1 => A3(38), B2 => 
                           n158, C1 => A2(38), C2 => n150, ZN => n244);
   U125 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U126 : AOI22_X1 port map( A1 => A0(39), A2 => n141, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U127 : AOI222_X1 port map( A1 => A1(39), A2 => n166, B1 => A3(39), B2 => 
                           n158, C1 => A2(39), C2 => n150, ZN => n246);
   U128 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U129 : AOI22_X1 port map( A1 => A0(47), A2 => n142, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U130 : AOI222_X1 port map( A1 => A1(47), A2 => n167, B1 => A3(47), B2 => 
                           n159, C1 => A2(47), C2 => n151, ZN => n264);
   U131 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U132 : AOI22_X1 port map( A1 => A0(40), A2 => n141, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U133 : AOI222_X1 port map( A1 => A1(40), A2 => n166, B1 => A3(40), B2 => 
                           n158, C1 => A2(40), C2 => n150, ZN => n250);
   U134 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U135 : AOI22_X1 port map( A1 => A0(41), A2 => n141, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U136 : AOI222_X1 port map( A1 => A1(41), A2 => n166, B1 => A3(41), B2 => 
                           n158, C1 => A2(41), C2 => n150, ZN => n252);
   U137 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U138 : AOI22_X1 port map( A1 => A0(42), A2 => n142, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U139 : AOI222_X1 port map( A1 => A1(42), A2 => n167, B1 => A3(42), B2 => 
                           n159, C1 => A2(42), C2 => n151, ZN => n254);
   U140 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U141 : AOI22_X1 port map( A1 => A0(48), A2 => n142, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U142 : AOI222_X1 port map( A1 => A1(48), A2 => n167, B1 => A3(48), B2 => 
                           n159, C1 => A2(48), C2 => n151, ZN => n266);
   U143 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U144 : AOI22_X1 port map( A1 => A0(43), A2 => n142, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U145 : AOI222_X1 port map( A1 => A1(43), A2 => n167, B1 => A3(43), B2 => 
                           n159, C1 => A2(43), C2 => n151, ZN => n256);
   U146 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U147 : AOI22_X1 port map( A1 => A0(44), A2 => n142, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U148 : AOI222_X1 port map( A1 => A1(44), A2 => n167, B1 => A3(44), B2 => 
                           n159, C1 => A2(44), C2 => n151, ZN => n258);
   U149 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U150 : AOI22_X1 port map( A1 => A0(49), A2 => n142, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U151 : AOI222_X1 port map( A1 => A1(49), A2 => n167, B1 => A3(49), B2 => 
                           n159, C1 => A2(49), C2 => n151, ZN => n268);
   U152 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U153 : AOI22_X1 port map( A1 => A0(45), A2 => n142, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U154 : AOI222_X1 port map( A1 => A1(45), A2 => n167, B1 => A3(45), B2 => 
                           n159, C1 => A2(45), C2 => n151, ZN => n260);
   U155 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U156 : AOI22_X1 port map( A1 => A0(50), A2 => n142, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U157 : AOI222_X1 port map( A1 => A1(50), A2 => n167, B1 => A3(50), B2 => 
                           n159, C1 => A2(50), C2 => n151, ZN => n272);
   U158 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U159 : AOI22_X1 port map( A1 => A0(51), A2 => n142, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U160 : AOI222_X1 port map( A1 => A1(51), A2 => n167, B1 => A3(51), B2 => 
                           n159, C1 => A2(51), C2 => n151, ZN => n274);
   U161 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U162 : AOI22_X1 port map( A1 => A0(52), A2 => n142, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U163 : AOI222_X1 port map( A1 => A1(52), A2 => n167, B1 => A3(52), B2 => 
                           n159, C1 => A2(52), C2 => n151, ZN => n276);
   U164 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U165 : AOI22_X1 port map( A1 => A0(53), A2 => n143, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U166 : AOI222_X1 port map( A1 => A1(53), A2 => n168, B1 => A3(53), B2 => 
                           n160, C1 => A2(53), C2 => n152, ZN => n278);
   U167 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U168 : AOI22_X1 port map( A1 => A0(54), A2 => n143, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U169 : AOI222_X1 port map( A1 => A1(54), A2 => n168, B1 => A3(54), B2 => 
                           n160, C1 => A2(54), C2 => n152, ZN => n280);
   U170 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U171 : AOI22_X1 port map( A1 => A0(55), A2 => n143, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U172 : AOI222_X1 port map( A1 => A1(55), A2 => n168, B1 => A3(55), B2 => 
                           n160, C1 => A2(55), C2 => n152, ZN => n282);
   U173 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U174 : AOI22_X1 port map( A1 => A0(56), A2 => n143, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U175 : AOI222_X1 port map( A1 => A1(56), A2 => n168, B1 => A3(56), B2 => 
                           n160, C1 => A2(56), C2 => n152, ZN => n284);
   U176 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U177 : AOI22_X1 port map( A1 => A0(57), A2 => n143, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U178 : AOI222_X1 port map( A1 => A1(57), A2 => n168, B1 => A3(57), B2 => 
                           n160, C1 => A2(57), C2 => n152, ZN => n286);
   U179 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U180 : AOI22_X1 port map( A1 => A0(58), A2 => n143, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U181 : AOI222_X1 port map( A1 => A1(58), A2 => n168, B1 => A3(58), B2 => 
                           n160, C1 => A2(58), C2 => n152, ZN => n288);
   U182 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U183 : AOI22_X1 port map( A1 => A0(59), A2 => n143, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U184 : AOI222_X1 port map( A1 => A1(59), A2 => n168, B1 => A3(59), B2 => 
                           n160, C1 => A2(59), C2 => n152, ZN => n290);
   U185 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U186 : AOI22_X1 port map( A1 => A0(60), A2 => n143, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U187 : AOI222_X1 port map( A1 => A1(60), A2 => n168, B1 => A3(60), B2 => 
                           n160, C1 => A2(60), C2 => n152, ZN => n294);
   U188 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U189 : AOI22_X1 port map( A1 => A0(61), A2 => n143, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U190 : AOI222_X1 port map( A1 => A1(61), A2 => n168, B1 => A3(61), B2 => 
                           n160, C1 => A2(61), C2 => n152, ZN => n296);
   U191 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U192 : AOI22_X1 port map( A1 => A0(62), A2 => n143, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U193 : AOI222_X1 port map( A1 => A1(62), A2 => n168, B1 => A3(62), B2 => 
                           n160, C1 => A2(62), C2 => n152, ZN => n298);
   U194 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U195 : AOI22_X1 port map( A1 => A0(63), A2 => n143, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U196 : AOI222_X1 port map( A1 => A1(63), A2 => n168, B1 => A3(63), B2 => 
                           n160, C1 => A2(63), C2 => n152, ZN => n300);
   U197 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U198 : AOI22_X1 port map( A1 => A0(0), A2 => n139, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U199 : AOI222_X1 port map( A1 => A1(0), A2 => n164, B1 => A3(0), B2 => n156,
                           C1 => A2(0), C2 => n148, ZN => n182);
   U200 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U201 : AOI22_X1 port map( A1 => A0(1), A2 => n139, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U202 : AOI222_X1 port map( A1 => A1(1), A2 => n164, B1 => A3(1), B2 => n156,
                           C1 => A2(1), C2 => n148, ZN => n204);
   U203 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U204 : AOI22_X1 port map( A1 => A0(2), A2 => n140, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U205 : AOI222_X1 port map( A1 => A1(2), A2 => n165, B1 => A3(2), B2 => n157,
                           C1 => A2(2), C2 => n149, ZN => n226);
   U206 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U207 : AOI22_X1 port map( A1 => A0(3), A2 => n141, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U208 : AOI222_X1 port map( A1 => A1(3), A2 => n166, B1 => A3(3), B2 => n158,
                           C1 => A2(3), C2 => n150, ZN => n248);
   U209 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U210 : AOI22_X1 port map( A1 => A0(4), A2 => n142, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U211 : AOI222_X1 port map( A1 => A1(4), A2 => n167, B1 => A3(4), B2 => n159,
                           C1 => A2(4), C2 => n151, ZN => n270);
   U212 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U213 : AOI22_X1 port map( A1 => A0(5), A2 => n143, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U214 : AOI222_X1 port map( A1 => A1(5), A2 => n168, B1 => A3(5), B2 => n160,
                           C1 => A2(5), C2 => n152, ZN => n292);
   U215 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U216 : AOI22_X1 port map( A1 => A0(6), A2 => n144, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U217 : AOI222_X1 port map( A1 => A1(6), A2 => n169, B1 => A3(6), B2 => n161,
                           C1 => A2(6), C2 => n153, ZN => n302);
   U218 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U219 : AOI22_X1 port map( A1 => A0(7), A2 => n144, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U220 : AOI222_X1 port map( A1 => A1(7), A2 => n169, B1 => A3(7), B2 => n161,
                           C1 => A2(7), C2 => n153, ZN => n304);
   U221 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U222 : AOI22_X1 port map( A1 => A0(8), A2 => n144, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U223 : AOI222_X1 port map( A1 => A1(8), A2 => n169, B1 => A3(8), B2 => n161,
                           C1 => A2(8), C2 => n153, ZN => n306);
   U224 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => O(9));
   U225 : AOI22_X1 port map( A1 => A0(9), A2 => n144, B1 => n178, B2 => A4(9), 
                           ZN => n310);
   U226 : AOI222_X1 port map( A1 => A1(9), A2 => n169, B1 => A3(9), B2 => n161,
                           C1 => A2(9), C2 => n153, ZN => n309);
   U227 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U228 : AOI22_X1 port map( A1 => A0(10), A2 => n139, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U229 : AOI222_X1 port map( A1 => A1(10), A2 => n164, B1 => A3(10), B2 => 
                           n156, C1 => A2(10), C2 => n148, ZN => n184);
   U230 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U231 : AOI22_X1 port map( A1 => A0(11), A2 => n139, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U232 : AOI222_X1 port map( A1 => A1(11), A2 => n164, B1 => A3(11), B2 => 
                           n156, C1 => A2(11), C2 => n148, ZN => n186);
   U233 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U234 : AOI22_X1 port map( A1 => A0(12), A2 => n139, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U235 : AOI222_X1 port map( A1 => A1(12), A2 => n164, B1 => A3(12), B2 => 
                           n156, C1 => A2(12), C2 => n148, ZN => n188);
   U236 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U237 : AOI22_X1 port map( A1 => A0(13), A2 => n139, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U238 : AOI222_X1 port map( A1 => A1(13), A2 => n164, B1 => A3(13), B2 => 
                           n156, C1 => A2(13), C2 => n148, ZN => n190);
   U239 : AOI22_X1 port map( A1 => A0(18), A2 => n139, B1 => A4(18), B2 => n177
                           , ZN => n201);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_8 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_8;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_8 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n136, Z => n154);
   U2 : BUF_X1 port map( A => n171, Z => n170);
   U3 : BUF_X1 port map( A => n137, Z => n162);
   U4 : BUF_X1 port map( A => n136, Z => n153);
   U5 : BUF_X1 port map( A => n171, Z => n169);
   U6 : BUF_X1 port map( A => n137, Z => n161);
   U7 : BUF_X1 port map( A => n146, Z => n145);
   U8 : BUF_X1 port map( A => n146, Z => n144);
   U9 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U10 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n147);
   U14 : BUF_X1 port map( A => n170, Z => n163);
   U15 : BUF_X1 port map( A => n162, Z => n155);
   U16 : BUF_X1 port map( A => n154, Z => n148);
   U17 : BUF_X1 port map( A => n170, Z => n164);
   U18 : BUF_X1 port map( A => n162, Z => n156);
   U19 : BUF_X1 port map( A => n170, Z => n165);
   U20 : BUF_X1 port map( A => n154, Z => n149);
   U21 : BUF_X1 port map( A => n162, Z => n157);
   U22 : BUF_X1 port map( A => n169, Z => n166);
   U23 : BUF_X1 port map( A => n153, Z => n150);
   U24 : BUF_X1 port map( A => n161, Z => n158);
   U25 : BUF_X1 port map( A => n169, Z => n167);
   U26 : BUF_X1 port map( A => n153, Z => n151);
   U27 : BUF_X1 port map( A => n161, Z => n159);
   U28 : BUF_X1 port map( A => n145, Z => n138);
   U29 : BUF_X1 port map( A => n145, Z => n140);
   U30 : BUF_X1 port map( A => n144, Z => n141);
   U31 : BUF_X1 port map( A => n144, Z => n142);
   U32 : BUF_X1 port map( A => n145, Z => n139);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n177);
   U38 : BUF_X1 port map( A => n179, Z => n176);
   U39 : BUF_X1 port map( A => n180, Z => n175);
   U40 : BUF_X1 port map( A => n180, Z => n174);
   U41 : BUF_X1 port map( A => n180, Z => n173);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U49 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177,
                           ZN => n197);
   U50 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => n155
                           , C1 => A2(16), C2 => n147, ZN => n196);
   U51 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U52 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177,
                           ZN => n199);
   U53 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U54 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U55 : BUF_X1 port map( A => sel(2), Z => n172);
   U56 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U57 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U58 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U59 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U60 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U61 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U62 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U63 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U64 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U65 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U66 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U67 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U68 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U69 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U70 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U71 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => n156
                           , C1 => A2(26), C2 => n148, ZN => n218);
   U72 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U73 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U74 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => n157
                           , C1 => A2(33), C2 => n149, ZN => n234);
   U75 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U76 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U77 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U78 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U79 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U80 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => n157
                           , C1 => A2(31), C2 => n149, ZN => n230);
   U81 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U82 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U83 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => n156
                           , C1 => A2(27), C2 => n148, ZN => n220);
   U84 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U85 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U86 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => n157
                           , C1 => A2(35), C2 => n149, ZN => n238);
   U87 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U88 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176,
                           ZN => n223);
   U89 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => n156
                           , C1 => A2(28), C2 => n148, ZN => n222);
   U90 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U91 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U92 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U93 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U94 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U95 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => n156
                           , C1 => A2(29), C2 => n148, ZN => n224);
   U96 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U97 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U98 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U99 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U100 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U101 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => 
                           n156, C1 => A2(30), C2 => n148, ZN => n228);
   U102 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U103 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => 
                           n157, C1 => A2(32), C2 => n149, ZN => n232);
   U104 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U105 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U106 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U107 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => 
                           n157, C1 => A2(38), C2 => n149, ZN => n244);
   U108 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U109 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U110 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => 
                           n157, C1 => A2(39), C2 => n149, ZN => n246);
   U111 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U112 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U113 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U114 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U115 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U116 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => 
                           n157, C1 => A2(40), C2 => n149, ZN => n250);
   U117 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U118 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U119 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => 
                           n157, C1 => A2(41), C2 => n149, ZN => n252);
   U120 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U121 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U122 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U123 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U124 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U125 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => 
                           n158, C1 => A2(42), C2 => n150, ZN => n254);
   U126 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U127 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U128 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => 
                           n158, C1 => A2(43), C2 => n150, ZN => n256);
   U129 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U130 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U131 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U132 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U133 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U134 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U135 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U136 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U137 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => 
                           n158, C1 => A2(45), C2 => n150, ZN => n260);
   U138 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U139 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U140 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U141 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U142 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U143 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U144 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U145 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U146 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => 
                           n158, C1 => A2(47), C2 => n150, ZN => n264);
   U147 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U148 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U149 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U150 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U151 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U152 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U153 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U154 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U155 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U156 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U157 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U158 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U159 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U160 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U161 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U162 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U163 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U164 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U165 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U166 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U167 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U168 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U169 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U170 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U171 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U172 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U173 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U174 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U175 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U176 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U177 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U178 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U179 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U180 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U181 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U182 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U183 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U184 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U185 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U186 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U187 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U188 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U189 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U190 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U191 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U192 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U193 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U194 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U195 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U196 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U197 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U198 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U199 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U200 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U201 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U202 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U203 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U204 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U205 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U206 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U207 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U208 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U209 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U210 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U211 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U212 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U213 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U214 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U215 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U216 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U217 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U218 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U219 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U220 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U221 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U222 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U223 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U224 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U225 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U226 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U227 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U228 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U229 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U230 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U231 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U232 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U233 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U234 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U235 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);
   U236 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U237 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U238 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U239 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U240 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_7 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_7;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n147);
   U14 : BUF_X1 port map( A => n170, Z => n163);
   U15 : BUF_X1 port map( A => n162, Z => n155);
   U16 : BUF_X1 port map( A => n170, Z => n164);
   U17 : BUF_X1 port map( A => n154, Z => n148);
   U18 : BUF_X1 port map( A => n162, Z => n156);
   U19 : BUF_X1 port map( A => n170, Z => n165);
   U20 : BUF_X1 port map( A => n154, Z => n149);
   U21 : BUF_X1 port map( A => n162, Z => n157);
   U22 : BUF_X1 port map( A => n169, Z => n166);
   U23 : BUF_X1 port map( A => n153, Z => n150);
   U24 : BUF_X1 port map( A => n161, Z => n158);
   U25 : BUF_X1 port map( A => n169, Z => n167);
   U26 : BUF_X1 port map( A => n153, Z => n151);
   U27 : BUF_X1 port map( A => n161, Z => n159);
   U28 : BUF_X1 port map( A => n145, Z => n138);
   U29 : BUF_X1 port map( A => n145, Z => n140);
   U30 : BUF_X1 port map( A => n144, Z => n141);
   U31 : BUF_X1 port map( A => n144, Z => n142);
   U32 : BUF_X1 port map( A => n145, Z => n139);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n177);
   U38 : BUF_X1 port map( A => n179, Z => n176);
   U39 : BUF_X1 port map( A => n180, Z => n175);
   U40 : BUF_X1 port map( A => n180, Z => n174);
   U41 : BUF_X1 port map( A => n180, Z => n173);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U49 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177,
                           ZN => n201);
   U50 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => n155
                           , C1 => A2(18), C2 => n147, ZN => n200);
   U51 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U52 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177,
                           ZN => n203);
   U53 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => n155
                           , C1 => A2(19), C2 => n147, ZN => n202);
   U54 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U55 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U56 : BUF_X1 port map( A => sel(2), Z => n172);
   U57 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U58 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U59 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => n156
                           , C1 => A2(21), C2 => n148, ZN => n208);
   U60 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U61 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U62 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U63 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => n156
                           , C1 => A2(23), C2 => n148, ZN => n212);
   U64 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U65 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => n156
                           , C1 => A2(24), C2 => n148, ZN => n214);
   U66 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U67 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U68 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => n156
                           , C1 => A2(25), C2 => n148, ZN => n216);
   U69 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U70 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => n156
                           , C1 => A2(26), C2 => n148, ZN => n218);
   U71 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U72 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U73 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => n156
                           , C1 => A2(27), C2 => n148, ZN => n220);
   U74 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U75 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => n156
                           , C1 => A2(28), C2 => n148, ZN => n222);
   U76 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U77 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U78 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => n157
                           , C1 => A2(35), C2 => n149, ZN => n238);
   U79 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U80 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U81 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => n156
                           , C1 => A2(29), C2 => n148, ZN => n224);
   U82 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U83 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U84 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U85 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U86 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U87 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => n157
                           , C1 => A2(33), C2 => n149, ZN => n234);
   U88 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U89 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U90 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U91 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U92 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176,
                           ZN => n229);
   U93 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => n156
                           , C1 => A2(30), C2 => n148, ZN => n228);
   U94 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U95 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U96 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U97 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U98 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U99 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => n157
                           , C1 => A2(31), C2 => n149, ZN => n230);
   U100 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U101 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175
                           , ZN => n247);
   U102 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => 
                           n157, C1 => A2(39), C2 => n149, ZN => n246);
   U103 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U104 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U105 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => 
                           n157, C1 => A2(32), C2 => n149, ZN => n232);
   U106 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U107 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U108 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => 
                           n157, C1 => A2(40), C2 => n149, ZN => n250);
   U109 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U110 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U111 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => 
                           n157, C1 => A2(41), C2 => n149, ZN => n252);
   U112 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U113 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U114 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U115 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U116 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U117 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => 
                           n157, C1 => A2(34), C2 => n149, ZN => n236);
   U118 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U119 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U120 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => 
                           n158, C1 => A2(42), C2 => n150, ZN => n254);
   U121 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U122 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U123 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => 
                           n158, C1 => A2(43), C2 => n150, ZN => n256);
   U124 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U125 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U126 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U127 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U128 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U129 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U130 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U131 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U132 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => 
                           n158, C1 => A2(45), C2 => n150, ZN => n260);
   U133 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U134 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U135 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U136 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U137 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U138 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U139 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U140 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U141 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => 
                           n158, C1 => A2(47), C2 => n150, ZN => n264);
   U142 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U143 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U144 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U145 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U146 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U147 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U148 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U149 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U150 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U151 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U152 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U153 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U154 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U155 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U156 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U157 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U158 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U159 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U160 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U161 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U162 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U163 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U164 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U165 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U166 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U167 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U168 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U169 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U170 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U171 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U172 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U173 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U174 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U175 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U176 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U177 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U178 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U179 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U180 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U181 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U182 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U183 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U184 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U185 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U186 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U187 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U188 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U189 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U190 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U191 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U192 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U193 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U194 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U195 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U196 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U197 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U198 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U199 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U200 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U201 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U202 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U203 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U204 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U205 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U206 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U207 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U208 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U209 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U210 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U211 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U212 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U213 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U214 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U215 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U216 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U217 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U218 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U219 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U220 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U221 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U222 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U223 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U224 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U225 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U226 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U227 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U228 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U229 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U230 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U231 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U232 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U233 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U234 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U235 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U236 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U237 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U238 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U239 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U240 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176
                           , ZN => n215);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_6 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_6;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_6 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n164);
   U15 : BUF_X1 port map( A => n162, Z => n156);
   U16 : BUF_X1 port map( A => n170, Z => n165);
   U17 : BUF_X1 port map( A => n154, Z => n149);
   U18 : BUF_X1 port map( A => n162, Z => n157);
   U19 : BUF_X1 port map( A => n169, Z => n166);
   U20 : BUF_X1 port map( A => n153, Z => n150);
   U21 : BUF_X1 port map( A => n161, Z => n158);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n153, Z => n151);
   U24 : BUF_X1 port map( A => n161, Z => n159);
   U25 : BUF_X1 port map( A => n145, Z => n138);
   U26 : BUF_X1 port map( A => n145, Z => n140);
   U27 : BUF_X1 port map( A => n144, Z => n141);
   U28 : BUF_X1 port map( A => n144, Z => n142);
   U29 : BUF_X1 port map( A => n162, Z => n155);
   U30 : BUF_X1 port map( A => n154, Z => n147);
   U31 : BUF_X1 port map( A => n170, Z => n163);
   U32 : BUF_X1 port map( A => n145, Z => n139);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n177);
   U38 : BUF_X1 port map( A => n179, Z => n176);
   U39 : BUF_X1 port map( A => n180, Z => n175);
   U40 : BUF_X1 port map( A => n180, Z => n174);
   U41 : BUF_X1 port map( A => n180, Z => n173);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U49 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177,
                           ZN => n207);
   U50 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => n156
                           , C1 => A2(20), C2 => n148, ZN => n206);
   U51 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U52 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177,
                           ZN => n209);
   U53 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => n156
                           , C1 => A2(21), C2 => n148, ZN => n208);
   U54 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U55 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U56 : BUF_X1 port map( A => sel(2), Z => n172);
   U57 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U58 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U59 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U60 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U61 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => n156
                           , C1 => A2(26), C2 => n148, ZN => n218);
   U62 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U63 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U64 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U65 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => n156
                           , C1 => A2(28), C2 => n148, ZN => n222);
   U66 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U67 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U68 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U69 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => n156
                           , C1 => A2(30), C2 => n148, ZN => n228);
   U70 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U71 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U72 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => n157
                           , C1 => A2(31), C2 => n149, ZN => n230);
   U73 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U74 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U75 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => n157
                           , C1 => A2(39), C2 => n149, ZN => n246);
   U76 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U77 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176,
                           ZN => n233);
   U78 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => n157
                           , C1 => A2(32), C2 => n149, ZN => n232);
   U79 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U80 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175,
                           ZN => n251);
   U81 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => n157
                           , C1 => A2(40), C2 => n149, ZN => n250);
   U82 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U83 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U84 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => n157
                           , C1 => A2(33), C2 => n149, ZN => n234);
   U85 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U86 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U87 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U88 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U89 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175,
                           ZN => n253);
   U90 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => n157
                           , C1 => A2(41), C2 => n149, ZN => n252);
   U91 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U92 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U93 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U94 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U95 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U96 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U97 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U98 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U99 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => n157
                           , C1 => A2(35), C2 => n149, ZN => n238);
   U100 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U101 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U102 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => 
                           n158, C1 => A2(42), C2 => n150, ZN => n254);
   U103 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U104 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U105 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => 
                           n158, C1 => A2(43), C2 => n150, ZN => n256);
   U106 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U107 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175
                           , ZN => n241);
   U108 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => 
                           n157, C1 => A2(36), C2 => n149, ZN => n240);
   U109 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U110 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U111 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U112 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U113 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U114 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U115 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U116 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U117 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => 
                           n158, C1 => A2(45), C2 => n150, ZN => n260);
   U118 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U119 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U120 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U121 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U122 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U123 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U124 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U125 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U126 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => 
                           n158, C1 => A2(47), C2 => n150, ZN => n264);
   U127 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U128 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U129 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U130 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U131 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U132 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U133 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U134 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U135 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U136 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U137 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U138 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U139 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U140 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U141 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U142 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U143 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U144 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U145 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U146 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U147 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U148 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U149 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U150 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U151 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U152 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U153 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U154 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U155 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U156 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U157 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U158 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U159 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U160 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U161 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U162 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U163 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U164 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U165 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U166 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U167 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U168 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U169 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U170 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U171 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U172 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U173 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U174 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U175 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U176 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U177 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U178 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U179 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U180 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U181 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U182 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U183 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U184 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U185 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U186 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U187 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U188 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U189 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U190 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U191 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U192 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U193 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U194 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U195 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U196 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U197 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U198 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U199 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U200 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U201 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U202 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U203 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U204 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U205 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U206 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U207 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U208 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U209 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U210 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U211 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U212 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U213 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U214 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U215 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U216 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U217 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U218 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U219 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U220 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U221 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U222 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U223 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U224 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U225 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U226 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U227 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U228 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U229 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U230 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);
   U231 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U232 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U233 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U234 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U235 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U236 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => 
                           n156, C1 => A2(27), C2 => n148, ZN => n220);
   U237 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U238 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U239 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U240 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_5 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_5;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n164);
   U15 : BUF_X1 port map( A => n162, Z => n156);
   U16 : BUF_X1 port map( A => n170, Z => n165);
   U17 : BUF_X1 port map( A => n154, Z => n149);
   U18 : BUF_X1 port map( A => n162, Z => n157);
   U19 : BUF_X1 port map( A => n169, Z => n166);
   U20 : BUF_X1 port map( A => n153, Z => n150);
   U21 : BUF_X1 port map( A => n161, Z => n158);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n153, Z => n151);
   U24 : BUF_X1 port map( A => n161, Z => n159);
   U25 : BUF_X1 port map( A => n145, Z => n138);
   U26 : BUF_X1 port map( A => n144, Z => n141);
   U27 : BUF_X1 port map( A => n144, Z => n142);
   U28 : BUF_X1 port map( A => n162, Z => n155);
   U29 : BUF_X1 port map( A => n145, Z => n140);
   U30 : BUF_X1 port map( A => n154, Z => n147);
   U31 : BUF_X1 port map( A => n170, Z => n163);
   U32 : BUF_X1 port map( A => n145, Z => n139);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n176);
   U38 : BUF_X1 port map( A => n180, Z => n175);
   U39 : BUF_X1 port map( A => n180, Z => n174);
   U40 : BUF_X1 port map( A => n180, Z => n173);
   U41 : BUF_X1 port map( A => n179, Z => n177);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U49 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177,
                           ZN => n211);
   U50 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => n156
                           , C1 => A2(22), C2 => n148, ZN => n210);
   U51 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U52 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176,
                           ZN => n213);
   U53 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U54 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U55 : BUF_X1 port map( A => sel(2), Z => n172);
   U56 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U57 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U58 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U59 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U60 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => n156
                           , C1 => A2(28), C2 => n148, ZN => n222);
   U61 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U62 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U63 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U64 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U65 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U66 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U67 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => n157
                           , C1 => A2(32), C2 => n149, ZN => n232);
   U68 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U69 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U70 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => n157
                           , C1 => A2(33), C2 => n149, ZN => n234);
   U71 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U72 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175,
                           ZN => n253);
   U73 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => n157
                           , C1 => A2(41), C2 => n149, ZN => n252);
   U74 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U75 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U76 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U77 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U78 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175,
                           ZN => n255);
   U79 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => n158
                           , C1 => A2(42), C2 => n150, ZN => n254);
   U80 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U81 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U82 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => n157
                           , C1 => A2(35), C2 => n149, ZN => n238);
   U83 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U84 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U85 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => n157
                           , C1 => A2(39), C2 => n149, ZN => n246);
   U86 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U87 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175,
                           ZN => n257);
   U88 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => n158
                           , C1 => A2(43), C2 => n150, ZN => n256);
   U89 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U90 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U91 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U92 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U93 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175,
                           ZN => n251);
   U94 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => n157
                           , C1 => A2(40), C2 => n149, ZN => n250);
   U95 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U96 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U97 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U98 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U99 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174,
                           ZN => n259);
   U100 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U101 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U102 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U103 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => 
                           n158, C1 => A2(45), C2 => n150, ZN => n260);
   U104 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U105 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175
                           , ZN => n245);
   U106 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => 
                           n157, C1 => A2(38), C2 => n149, ZN => n244);
   U107 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U108 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U109 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U110 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U111 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U112 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U113 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U114 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U115 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => 
                           n158, C1 => A2(47), C2 => n150, ZN => n264);
   U116 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U117 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U118 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U119 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U120 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U121 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U122 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U123 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U124 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U125 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U126 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U127 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U128 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U129 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U130 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U131 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U132 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U133 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U134 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U135 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U136 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U137 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U138 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U139 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U140 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U141 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U142 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U143 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U144 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U145 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U146 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U147 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U148 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U149 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U150 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U151 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U152 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U153 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U154 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U155 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U156 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U157 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U158 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U159 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U160 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U161 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U162 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U163 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U164 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U165 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U166 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U167 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U168 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U169 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U170 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U171 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U172 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U173 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U174 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U175 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U176 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U177 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U178 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U179 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U180 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U181 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U182 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U183 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U184 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U185 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U186 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U187 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U188 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U189 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U190 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U191 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U192 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U193 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U194 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U195 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U196 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U197 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U198 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U199 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U200 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U201 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U202 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U203 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U204 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U205 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U206 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U207 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U208 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U209 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U210 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U211 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U212 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U213 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U214 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U215 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U216 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U217 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U218 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U219 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U220 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U221 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U222 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U223 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U224 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U225 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U226 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U227 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U228 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U229 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => 
                           n157, C1 => A2(31), C2 => n149, ZN => n230);
   U230 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U231 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => 
                           n156, C1 => A2(30), C2 => n148, ZN => n228);
   U232 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => 
                           n156, C1 => A2(26), C2 => n148, ZN => n218);
   U233 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U234 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U235 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);
   U236 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U237 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U238 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);
   U239 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U240 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => 
                           n156, C1 => A2(27), C2 => n148, ZN => n220);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_4 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_4;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n164);
   U15 : BUF_X1 port map( A => n162, Z => n156);
   U16 : BUF_X1 port map( A => n170, Z => n165);
   U17 : BUF_X1 port map( A => n154, Z => n149);
   U18 : BUF_X1 port map( A => n162, Z => n157);
   U19 : BUF_X1 port map( A => n169, Z => n166);
   U20 : BUF_X1 port map( A => n153, Z => n150);
   U21 : BUF_X1 port map( A => n161, Z => n158);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n153, Z => n151);
   U24 : BUF_X1 port map( A => n161, Z => n159);
   U25 : BUF_X1 port map( A => n145, Z => n138);
   U26 : BUF_X1 port map( A => n144, Z => n141);
   U27 : BUF_X1 port map( A => n144, Z => n142);
   U28 : BUF_X1 port map( A => n162, Z => n155);
   U29 : BUF_X1 port map( A => n154, Z => n147);
   U30 : BUF_X1 port map( A => n170, Z => n163);
   U31 : BUF_X1 port map( A => n145, Z => n140);
   U32 : BUF_X1 port map( A => n145, Z => n139);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n176);
   U38 : BUF_X1 port map( A => n180, Z => n175);
   U39 : BUF_X1 port map( A => n180, Z => n174);
   U40 : BUF_X1 port map( A => n180, Z => n173);
   U41 : BUF_X1 port map( A => n179, Z => n177);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U49 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176,
                           ZN => n215);
   U50 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => n156
                           , C1 => A2(24), C2 => n148, ZN => n214);
   U51 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U52 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176,
                           ZN => n217);
   U53 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => n156
                           , C1 => A2(25), C2 => n148, ZN => n216);
   U54 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U55 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U56 : BUF_X1 port map( A => sel(2), Z => n172);
   U57 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U58 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U59 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U60 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U61 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => n156
                           , C1 => A2(30), C2 => n148, ZN => n228);
   U62 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U63 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U64 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U65 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => n157
                           , C1 => A2(32), C2 => n149, ZN => n232);
   U66 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U67 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U68 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U69 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U70 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U71 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U72 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => n157
                           , C1 => A2(35), C2 => n149, ZN => n238);
   U73 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U74 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175,
                           ZN => n257);
   U75 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => n158
                           , C1 => A2(43), C2 => n150, ZN => n256);
   U76 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U77 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U78 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U79 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U80 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174,
                           ZN => n259);
   U81 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => n158
                           , C1 => A2(44), C2 => n150, ZN => n258);
   U82 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U83 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U84 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U85 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U86 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175,
                           ZN => n253);
   U87 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => n157
                           , C1 => A2(41), C2 => n149, ZN => n252);
   U88 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U89 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174,
                           ZN => n261);
   U90 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => n158
                           , C1 => A2(45), C2 => n150, ZN => n260);
   U91 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U92 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U93 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U94 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U95 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175,
                           ZN => n255);
   U96 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => n158
                           , C1 => A2(42), C2 => n150, ZN => n254);
   U97 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U98 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U99 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => n157
                           , C1 => A2(39), C2 => n149, ZN => n246);
   U100 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U101 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U102 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U103 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U104 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174
                           , ZN => n265);
   U105 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => 
                           n158, C1 => A2(47), C2 => n150, ZN => n264);
   U106 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U107 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U108 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => 
                           n157, C1 => A2(40), C2 => n149, ZN => n250);
   U109 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U110 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U111 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U112 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U113 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U114 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U115 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U116 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U117 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U118 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U119 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U120 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U121 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U122 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U123 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U124 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U125 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U126 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U127 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U128 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U129 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U130 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U131 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U132 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U133 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U134 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U135 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U136 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U137 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U138 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U139 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U140 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U141 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U142 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U143 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U144 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U145 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U146 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U147 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U148 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U149 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U150 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U151 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U152 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U153 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U154 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U155 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U156 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U157 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U158 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U159 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U160 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U161 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U162 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U163 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U164 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U165 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U166 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U167 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U168 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U169 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U170 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U171 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U172 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U173 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U174 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U175 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U176 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U177 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U178 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U179 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U180 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U181 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U182 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U183 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U184 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U185 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U186 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U187 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U188 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U189 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U190 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U191 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U192 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U193 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U194 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U195 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U196 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U197 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U198 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U199 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U200 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U201 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U202 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U203 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U204 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U205 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U206 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U207 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U208 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U209 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U210 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U211 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U212 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U213 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U214 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U215 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U216 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U217 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U218 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U219 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U220 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U221 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U222 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U223 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U224 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U225 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U226 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U227 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U228 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U229 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U230 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => 
                           n157, C1 => A2(33), C2 => n149, ZN => n234);
   U231 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U232 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => 
                           n156, C1 => A2(26), C2 => n148, ZN => n218);
   U233 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => 
                           n156, C1 => A2(28), C2 => n148, ZN => n222);
   U234 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176
                           , ZN => n225);
   U235 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U236 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => 
                           n157, C1 => A2(31), C2 => n149, ZN => n230);
   U237 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U238 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => 
                           n156, C1 => A2(27), C2 => n148, ZN => n220);
   U239 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U240 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_3 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_3;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n164);
   U15 : BUF_X1 port map( A => n162, Z => n156);
   U16 : BUF_X1 port map( A => n170, Z => n165);
   U17 : BUF_X1 port map( A => n154, Z => n149);
   U18 : BUF_X1 port map( A => n162, Z => n157);
   U19 : BUF_X1 port map( A => n169, Z => n166);
   U20 : BUF_X1 port map( A => n153, Z => n150);
   U21 : BUF_X1 port map( A => n161, Z => n158);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n153, Z => n151);
   U24 : BUF_X1 port map( A => n161, Z => n159);
   U25 : BUF_X1 port map( A => n145, Z => n138);
   U26 : BUF_X1 port map( A => n145, Z => n140);
   U27 : BUF_X1 port map( A => n144, Z => n141);
   U28 : BUF_X1 port map( A => n144, Z => n142);
   U29 : BUF_X1 port map( A => n162, Z => n155);
   U30 : BUF_X1 port map( A => n145, Z => n139);
   U31 : BUF_X1 port map( A => n154, Z => n147);
   U32 : BUF_X1 port map( A => n170, Z => n163);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n176);
   U38 : BUF_X1 port map( A => n180, Z => n175);
   U39 : BUF_X1 port map( A => n180, Z => n174);
   U40 : BUF_X1 port map( A => n180, Z => n173);
   U41 : BUF_X1 port map( A => n179, Z => n177);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U49 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176,
                           ZN => n219);
   U50 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => n156
                           , C1 => A2(26), C2 => n148, ZN => n218);
   U51 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U52 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176,
                           ZN => n221);
   U53 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => n156
                           , C1 => A2(27), C2 => n148, ZN => n220);
   U54 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U55 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176,
                           ZN => n223);
   U56 : BUF_X1 port map( A => sel(2), Z => n172);
   U57 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U58 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U59 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U60 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U61 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U62 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U63 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176,
                           ZN => n233);
   U64 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => n157
                           , C1 => A2(32), C2 => n149, ZN => n232);
   U65 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U66 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U67 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U68 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U69 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U70 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U71 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U72 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U73 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U74 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U75 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U76 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U77 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => n157
                           , C1 => A2(37), C2 => n149, ZN => n242);
   U78 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U79 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174,
                           ZN => n261);
   U80 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => n158
                           , C1 => A2(45), C2 => n150, ZN => n260);
   U81 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U82 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U83 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U84 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U85 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174,
                           ZN => n263);
   U86 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => n158
                           , C1 => A2(46), C2 => n150, ZN => n262);
   U87 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U88 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U89 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => n157
                           , C1 => A2(39), C2 => n149, ZN => n246);
   U90 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U91 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => n158
                           , C1 => A2(44), C2 => n150, ZN => n258);
   U92 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174,
                           ZN => n259);
   U93 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U94 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175,
                           ZN => n257);
   U95 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => n158
                           , C1 => A2(43), C2 => n150, ZN => n256);
   U96 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U97 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174,
                           ZN => n265);
   U98 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => n158
                           , C1 => A2(47), C2 => n150, ZN => n264);
   U99 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U100 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175
                           , ZN => n251);
   U101 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => 
                           n157, C1 => A2(40), C2 => n149, ZN => n250);
   U102 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U103 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175
                           , ZN => n253);
   U104 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => 
                           n157, C1 => A2(41), C2 => n149, ZN => n252);
   U105 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U106 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => 
                           n158, C1 => A2(42), C2 => n150, ZN => n254);
   U107 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175
                           , ZN => n255);
   U108 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U109 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174
                           , ZN => n267);
   U110 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => 
                           n158, C1 => A2(48), C2 => n150, ZN => n266);
   U111 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U112 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174
                           , ZN => n269);
   U113 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => 
                           n158, C1 => A2(49), C2 => n150, ZN => n268);
   U114 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U115 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U116 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U117 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U118 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U119 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U120 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U121 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U122 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U123 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U124 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U125 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U126 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U127 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U128 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U129 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U130 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U131 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U132 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U133 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U134 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U135 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U136 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U137 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U138 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U139 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U140 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U141 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U142 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U143 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U144 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U145 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U146 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U147 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U148 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U149 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U150 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U151 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U152 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U153 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U154 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U155 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U156 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U157 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U158 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U159 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U160 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U161 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U162 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U163 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U164 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U165 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U166 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U167 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U168 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U169 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U170 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U171 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U172 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U173 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U174 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U175 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U176 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U177 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U178 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U179 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U180 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U181 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U182 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U183 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U184 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U185 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U186 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U187 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U188 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U189 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U190 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U191 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U192 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U193 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U194 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U195 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U196 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U197 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U198 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U199 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U200 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U201 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U202 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U203 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U204 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U205 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U206 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U207 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U208 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U209 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U210 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U211 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U212 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U213 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U214 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U215 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U216 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U217 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U218 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U219 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U220 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U221 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U222 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U223 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U224 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U225 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U226 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U227 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U228 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U229 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U230 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U231 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U232 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U233 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);
   U234 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => 
                           n157, C1 => A2(35), C2 => n149, ZN => n238);
   U235 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => 
                           n156, C1 => A2(28), C2 => n148, ZN => n222);
   U236 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176
                           , ZN => n229);
   U237 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => 
                           n156, C1 => A2(30), C2 => n148, ZN => n228);
   U238 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => 
                           n157, C1 => A2(33), C2 => n149, ZN => n234);
   U239 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);
   U240 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => 
                           n157, C1 => A2(31), C2 => n149, ZN => n230);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_2 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_2;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n164);
   U15 : BUF_X1 port map( A => n162, Z => n156);
   U16 : BUF_X1 port map( A => n170, Z => n165);
   U17 : BUF_X1 port map( A => n154, Z => n149);
   U18 : BUF_X1 port map( A => n162, Z => n157);
   U19 : BUF_X1 port map( A => n169, Z => n166);
   U20 : BUF_X1 port map( A => n153, Z => n150);
   U21 : BUF_X1 port map( A => n161, Z => n158);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n153, Z => n151);
   U24 : BUF_X1 port map( A => n161, Z => n159);
   U25 : BUF_X1 port map( A => n145, Z => n138);
   U26 : BUF_X1 port map( A => n145, Z => n139);
   U27 : BUF_X1 port map( A => n144, Z => n141);
   U28 : BUF_X1 port map( A => n144, Z => n142);
   U29 : BUF_X1 port map( A => n162, Z => n155);
   U30 : BUF_X1 port map( A => n145, Z => n140);
   U31 : BUF_X1 port map( A => n154, Z => n147);
   U32 : BUF_X1 port map( A => n170, Z => n163);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n176);
   U38 : BUF_X1 port map( A => n180, Z => n175);
   U39 : BUF_X1 port map( A => n180, Z => n174);
   U40 : BUF_X1 port map( A => n180, Z => n173);
   U41 : BUF_X1 port map( A => n179, Z => n177);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U49 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176,
                           ZN => n223);
   U50 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => n156
                           , C1 => A2(28), C2 => n148, ZN => n222);
   U51 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U52 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176,
                           ZN => n225);
   U53 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U54 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176,
                           ZN => n229);
   U55 : BUF_X1 port map( A => sel(2), Z => n172);
   U56 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U57 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U58 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U59 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U60 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U61 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U62 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175,
                           ZN => n237);
   U63 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => n157
                           , C1 => A2(34), C2 => n149, ZN => n236);
   U64 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U65 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U66 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U67 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U68 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U69 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U70 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U71 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U72 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U73 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U74 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U75 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U76 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => n157
                           , C1 => A2(39), C2 => n149, ZN => n246);
   U77 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U78 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174,
                           ZN => n265);
   U79 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => n158
                           , C1 => A2(47), C2 => n150, ZN => n264);
   U80 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U81 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175,
                           ZN => n251);
   U82 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => n157
                           , C1 => A2(40), C2 => n149, ZN => n250);
   U83 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U84 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174,
                           ZN => n267);
   U85 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => n158
                           , C1 => A2(48), C2 => n150, ZN => n266);
   U86 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U87 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => n158
                           , C1 => A2(46), C2 => n150, ZN => n262);
   U88 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174,
                           ZN => n263);
   U89 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U90 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175,
                           ZN => n253);
   U91 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => n157
                           , C1 => A2(41), C2 => n149, ZN => n252);
   U92 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U93 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174,
                           ZN => n261);
   U94 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => n158
                           , C1 => A2(45), C2 => n150, ZN => n260);
   U95 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U96 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174,
                           ZN => n269);
   U97 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => n158
                           , C1 => A2(49), C2 => n150, ZN => n268);
   U98 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U99 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175,
                           ZN => n255);
   U100 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => 
                           n158, C1 => A2(42), C2 => n150, ZN => n254);
   U101 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U102 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175
                           , ZN => n257);
   U103 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => 
                           n158, C1 => A2(43), C2 => n150, ZN => n256);
   U104 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U105 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U106 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U107 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U108 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174
                           , ZN => n273);
   U109 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => 
                           n158, C1 => A2(50), C2 => n150, ZN => n272);
   U110 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U111 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174
                           , ZN => n275);
   U112 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => 
                           n158, C1 => A2(51), C2 => n150, ZN => n274);
   U113 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U114 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U115 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U116 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U117 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U118 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U119 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U120 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U121 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U122 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U123 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U124 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U125 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U126 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U127 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U128 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U129 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U130 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U131 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U132 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U133 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U134 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U135 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U136 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U137 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U138 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U139 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U140 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U141 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U142 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U143 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U144 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U145 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U146 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U147 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U148 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U149 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U150 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U151 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U152 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U153 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U154 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U155 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U156 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U157 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U158 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U159 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U160 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U161 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U162 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U163 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U164 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U165 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U166 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U167 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U168 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U169 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U170 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U171 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U172 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U173 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U174 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U175 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U176 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U177 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U178 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U179 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U180 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U181 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U182 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U183 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U184 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U185 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U186 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U187 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U188 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U189 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U190 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U191 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U192 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U193 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U194 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U195 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U196 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U197 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U198 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U199 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U200 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U201 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U202 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U203 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U204 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U205 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U206 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U207 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U208 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U209 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U210 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U211 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U212 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U213 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U214 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U215 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U216 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U217 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U218 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U219 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U220 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U221 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U222 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U223 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U224 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U225 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U226 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);
   U227 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U228 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U229 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => 
                           n156, C1 => A2(26), C2 => n148, ZN => n218);
   U230 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U231 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U232 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => 
                           n156, C1 => A2(27), C2 => n148, ZN => n220);
   U233 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);
   U234 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => 
                           n157, C1 => A2(37), C2 => n149, ZN => n242);
   U235 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176
                           , ZN => n233);
   U236 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => 
                           n157, C1 => A2(32), C2 => n149, ZN => n232);
   U237 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => 
                           n157, C1 => A2(35), C2 => n149, ZN => n238);
   U238 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => 
                           n156, C1 => A2(30), C2 => n148, ZN => n228);
   U239 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => 
                           n157, C1 => A2(31), C2 => n149, ZN => n230);
   U240 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => 
                           n157, C1 => A2(33), C2 => n149, ZN => n234);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_1 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_1;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => sel(1), A2 => n181, ZN => n136);
   U2 : AND2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n137);
   U3 : BUF_X1 port map( A => n136, Z => n154);
   U4 : BUF_X1 port map( A => n171, Z => n170);
   U5 : BUF_X1 port map( A => n137, Z => n162);
   U6 : BUF_X1 port map( A => n136, Z => n153);
   U7 : BUF_X1 port map( A => n171, Z => n169);
   U8 : BUF_X1 port map( A => n137, Z => n161);
   U9 : BUF_X1 port map( A => n146, Z => n145);
   U10 : BUF_X1 port map( A => n146, Z => n144);
   U11 : BUF_X1 port map( A => n172, Z => n179);
   U12 : BUF_X1 port map( A => n172, Z => n180);
   U13 : BUF_X1 port map( A => n154, Z => n148);
   U14 : BUF_X1 port map( A => n170, Z => n165);
   U15 : BUF_X1 port map( A => n154, Z => n149);
   U16 : BUF_X1 port map( A => n170, Z => n164);
   U17 : BUF_X1 port map( A => n162, Z => n157);
   U18 : BUF_X1 port map( A => n169, Z => n166);
   U19 : BUF_X1 port map( A => n153, Z => n150);
   U20 : BUF_X1 port map( A => n161, Z => n158);
   U21 : BUF_X1 port map( A => n153, Z => n151);
   U22 : BUF_X1 port map( A => n169, Z => n167);
   U23 : BUF_X1 port map( A => n161, Z => n159);
   U24 : BUF_X1 port map( A => n145, Z => n138);
   U25 : BUF_X1 port map( A => n145, Z => n139);
   U26 : BUF_X1 port map( A => n144, Z => n141);
   U27 : BUF_X1 port map( A => n144, Z => n142);
   U28 : BUF_X1 port map( A => n162, Z => n155);
   U29 : BUF_X1 port map( A => n162, Z => n156);
   U30 : BUF_X1 port map( A => n145, Z => n140);
   U31 : BUF_X1 port map( A => n154, Z => n147);
   U32 : BUF_X1 port map( A => n170, Z => n163);
   U33 : BUF_X1 port map( A => n144, Z => n143);
   U34 : BUF_X1 port map( A => n161, Z => n160);
   U35 : BUF_X1 port map( A => n153, Z => n152);
   U36 : BUF_X1 port map( A => n169, Z => n168);
   U37 : BUF_X1 port map( A => n179, Z => n176);
   U38 : BUF_X1 port map( A => n180, Z => n175);
   U39 : BUF_X1 port map( A => n180, Z => n174);
   U40 : BUF_X1 port map( A => n180, Z => n173);
   U41 : BUF_X1 port map( A => n179, Z => n177);
   U42 : BUF_X1 port map( A => n179, Z => n178);
   U43 : INV_X1 port map( A => sel(0), ZN => n181);
   U44 : BUF_X1 port map( A => n309, Z => n171);
   U45 : NOR2_X1 port map( A1 => n181, A2 => sel(1), ZN => n309);
   U46 : BUF_X1 port map( A => n308, Z => n146);
   U47 : NOR3_X1 port map( A1 => sel(1), A2 => n178, A3 => sel(0), ZN => n308);
   U48 : NAND2_X1 port map( A1 => n229, A2 => n228, ZN => O(30));
   U49 : AOI22_X1 port map( A1 => A0(30), A2 => n139, B1 => A4(30), B2 => n176,
                           ZN => n229);
   U50 : AOI222_X1 port map( A1 => A1(30), A2 => n164, B1 => A3(30), B2 => n156
                           , C1 => A2(30), C2 => n148, ZN => n228);
   U51 : NAND2_X1 port map( A1 => n231, A2 => n230, ZN => O(31));
   U52 : AOI22_X1 port map( A1 => A0(31), A2 => n140, B1 => A4(31), B2 => n176,
                           ZN => n231);
   U53 : AOI222_X1 port map( A1 => A1(31), A2 => n165, B1 => A3(31), B2 => n157
                           , C1 => A2(31), C2 => n149, ZN => n230);
   U54 : NAND2_X1 port map( A1 => n233, A2 => n232, ZN => O(32));
   U55 : AOI22_X1 port map( A1 => A0(32), A2 => n140, B1 => A4(32), B2 => n176,
                           ZN => n233);
   U56 : BUF_X1 port map( A => sel(2), Z => n172);
   U57 : NAND2_X1 port map( A1 => n235, A2 => n234, ZN => O(33));
   U58 : AOI22_X1 port map( A1 => A0(33), A2 => n140, B1 => A4(33), B2 => n176,
                           ZN => n235);
   U59 : NAND2_X1 port map( A1 => n237, A2 => n236, ZN => O(34));
   U60 : NAND2_X1 port map( A1 => n239, A2 => n238, ZN => O(35));
   U61 : AOI22_X1 port map( A1 => A0(35), A2 => n140, B1 => A4(35), B2 => n175,
                           ZN => n239);
   U62 : NAND2_X1 port map( A1 => n241, A2 => n240, ZN => O(36));
   U63 : AOI22_X1 port map( A1 => A0(36), A2 => n140, B1 => A4(36), B2 => n175,
                           ZN => n241);
   U64 : AOI222_X1 port map( A1 => A1(36), A2 => n165, B1 => A3(36), B2 => n157
                           , C1 => A2(36), C2 => n149, ZN => n240);
   U65 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => O(37));
   U66 : AOI22_X1 port map( A1 => A0(37), A2 => n140, B1 => A4(37), B2 => n175,
                           ZN => n243);
   U67 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => O(38));
   U68 : AOI22_X1 port map( A1 => A0(38), A2 => n140, B1 => A4(38), B2 => n175,
                           ZN => n245);
   U69 : AOI222_X1 port map( A1 => A1(38), A2 => n165, B1 => A3(38), B2 => n157
                           , C1 => A2(38), C2 => n149, ZN => n244);
   U70 : NAND2_X1 port map( A1 => n247, A2 => n246, ZN => O(39));
   U71 : AOI22_X1 port map( A1 => A0(39), A2 => n140, B1 => A4(39), B2 => n175,
                           ZN => n247);
   U72 : NAND2_X1 port map( A1 => n251, A2 => n250, ZN => O(40));
   U73 : AOI22_X1 port map( A1 => A0(40), A2 => n140, B1 => A4(40), B2 => n175,
                           ZN => n251);
   U74 : AOI222_X1 port map( A1 => A1(40), A2 => n165, B1 => A3(40), B2 => n157
                           , C1 => A2(40), C2 => n149, ZN => n250);
   U75 : NAND2_X1 port map( A1 => n253, A2 => n252, ZN => O(41));
   U76 : AOI22_X1 port map( A1 => A0(41), A2 => n140, B1 => A4(41), B2 => n175,
                           ZN => n253);
   U77 : AOI222_X1 port map( A1 => A1(41), A2 => n165, B1 => A3(41), B2 => n157
                           , C1 => A2(41), C2 => n149, ZN => n252);
   U78 : NAND2_X1 port map( A1 => n269, A2 => n268, ZN => O(49));
   U79 : AOI22_X1 port map( A1 => A0(49), A2 => n141, B1 => A4(49), B2 => n174,
                           ZN => n269);
   U80 : AOI222_X1 port map( A1 => A1(49), A2 => n166, B1 => A3(49), B2 => n158
                           , C1 => A2(49), C2 => n150, ZN => n268);
   U81 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => O(42));
   U82 : AOI22_X1 port map( A1 => A0(42), A2 => n141, B1 => A4(42), B2 => n175,
                           ZN => n255);
   U83 : AOI222_X1 port map( A1 => A1(42), A2 => n166, B1 => A3(42), B2 => n158
                           , C1 => A2(42), C2 => n150, ZN => n254);
   U84 : NAND2_X1 port map( A1 => n273, A2 => n272, ZN => O(50));
   U85 : AOI22_X1 port map( A1 => A0(50), A2 => n141, B1 => A4(50), B2 => n174,
                           ZN => n273);
   U86 : AOI222_X1 port map( A1 => A1(50), A2 => n166, B1 => A3(50), B2 => n158
                           , C1 => A2(50), C2 => n150, ZN => n272);
   U87 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => O(43));
   U88 : AOI22_X1 port map( A1 => A0(43), A2 => n141, B1 => A4(43), B2 => n175,
                           ZN => n257);
   U89 : AOI222_X1 port map( A1 => A1(43), A2 => n166, B1 => A3(43), B2 => n158
                           , C1 => A2(43), C2 => n150, ZN => n256);
   U90 : NAND2_X1 port map( A1 => n267, A2 => n266, ZN => O(48));
   U91 : AOI222_X1 port map( A1 => A1(48), A2 => n166, B1 => A3(48), B2 => n158
                           , C1 => A2(48), C2 => n150, ZN => n266);
   U92 : AOI22_X1 port map( A1 => A0(48), A2 => n141, B1 => A4(48), B2 => n174,
                           ZN => n267);
   U93 : NAND2_X1 port map( A1 => n265, A2 => n264, ZN => O(47));
   U94 : AOI22_X1 port map( A1 => A0(47), A2 => n141, B1 => A4(47), B2 => n174,
                           ZN => n265);
   U95 : AOI222_X1 port map( A1 => A1(47), A2 => n166, B1 => A3(47), B2 => n158
                           , C1 => A2(47), C2 => n150, ZN => n264);
   U96 : NAND2_X1 port map( A1 => n275, A2 => n274, ZN => O(51));
   U97 : AOI22_X1 port map( A1 => A0(51), A2 => n141, B1 => A4(51), B2 => n174,
                           ZN => n275);
   U98 : AOI222_X1 port map( A1 => A1(51), A2 => n166, B1 => A3(51), B2 => n158
                           , C1 => A2(51), C2 => n150, ZN => n274);
   U99 : NAND2_X1 port map( A1 => n259, A2 => n258, ZN => O(44));
   U100 : AOI22_X1 port map( A1 => A0(44), A2 => n141, B1 => A4(44), B2 => n174
                           , ZN => n259);
   U101 : AOI222_X1 port map( A1 => A1(44), A2 => n166, B1 => A3(44), B2 => 
                           n158, C1 => A2(44), C2 => n150, ZN => n258);
   U102 : NAND2_X1 port map( A1 => n261, A2 => n260, ZN => O(45));
   U103 : AOI22_X1 port map( A1 => A0(45), A2 => n141, B1 => A4(45), B2 => n174
                           , ZN => n261);
   U104 : AOI222_X1 port map( A1 => A1(45), A2 => n166, B1 => A3(45), B2 => 
                           n158, C1 => A2(45), C2 => n150, ZN => n260);
   U105 : NAND2_X1 port map( A1 => n263, A2 => n262, ZN => O(46));
   U106 : AOI222_X1 port map( A1 => A1(46), A2 => n166, B1 => A3(46), B2 => 
                           n158, C1 => A2(46), C2 => n150, ZN => n262);
   U107 : AOI22_X1 port map( A1 => A0(46), A2 => n141, B1 => A4(46), B2 => n174
                           , ZN => n263);
   U108 : NAND2_X1 port map( A1 => n277, A2 => n276, ZN => O(52));
   U109 : AOI22_X1 port map( A1 => A0(52), A2 => n141, B1 => A4(52), B2 => n175
                           , ZN => n277);
   U110 : AOI222_X1 port map( A1 => A1(52), A2 => n166, B1 => A3(52), B2 => 
                           n158, C1 => A2(52), C2 => n150, ZN => n276);
   U111 : NAND2_X1 port map( A1 => n279, A2 => n278, ZN => O(53));
   U112 : AOI22_X1 port map( A1 => A0(53), A2 => n142, B1 => A4(53), B2 => n174
                           , ZN => n279);
   U113 : AOI222_X1 port map( A1 => A1(53), A2 => n167, B1 => A3(53), B2 => 
                           n159, C1 => A2(53), C2 => n151, ZN => n278);
   U114 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => O(62));
   U115 : AOI22_X1 port map( A1 => A0(62), A2 => n142, B1 => A4(62), B2 => n173
                           , ZN => n299);
   U116 : AOI222_X1 port map( A1 => A1(62), A2 => n167, B1 => A3(62), B2 => 
                           n159, C1 => A2(62), C2 => n151, ZN => n298);
   U117 : NAND2_X1 port map( A1 => n281, A2 => n280, ZN => O(54));
   U118 : AOI22_X1 port map( A1 => A0(54), A2 => n142, B1 => A4(54), B2 => n174
                           , ZN => n281);
   U119 : AOI222_X1 port map( A1 => A1(54), A2 => n167, B1 => A3(54), B2 => 
                           n159, C1 => A2(54), C2 => n151, ZN => n280);
   U120 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => O(55));
   U121 : AOI22_X1 port map( A1 => A0(55), A2 => n142, B1 => A4(55), B2 => n174
                           , ZN => n283);
   U122 : AOI222_X1 port map( A1 => A1(55), A2 => n167, B1 => A3(55), B2 => 
                           n159, C1 => A2(55), C2 => n151, ZN => n282);
   U123 : NAND2_X1 port map( A1 => n301, A2 => n300, ZN => O(63));
   U124 : AOI22_X1 port map( A1 => A0(63), A2 => n142, B1 => A4(63), B2 => n173
                           , ZN => n301);
   U125 : AOI222_X1 port map( A1 => A1(63), A2 => n167, B1 => A3(63), B2 => 
                           n159, C1 => A2(63), C2 => n151, ZN => n300);
   U126 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => O(56));
   U127 : AOI22_X1 port map( A1 => A0(56), A2 => n142, B1 => A4(56), B2 => n173
                           , ZN => n285);
   U128 : AOI222_X1 port map( A1 => A1(56), A2 => n167, B1 => A3(56), B2 => 
                           n159, C1 => A2(56), C2 => n151, ZN => n284);
   U129 : NAND2_X1 port map( A1 => n287, A2 => n286, ZN => O(57));
   U130 : AOI22_X1 port map( A1 => A0(57), A2 => n142, B1 => A4(57), B2 => n173
                           , ZN => n287);
   U131 : AOI222_X1 port map( A1 => A1(57), A2 => n167, B1 => A3(57), B2 => 
                           n159, C1 => A2(57), C2 => n151, ZN => n286);
   U132 : NAND2_X1 port map( A1 => n289, A2 => n288, ZN => O(58));
   U133 : AOI22_X1 port map( A1 => A0(58), A2 => n142, B1 => A4(58), B2 => n173
                           , ZN => n289);
   U134 : AOI222_X1 port map( A1 => A1(58), A2 => n167, B1 => A3(58), B2 => 
                           n159, C1 => A2(58), C2 => n151, ZN => n288);
   U135 : NAND2_X1 port map( A1 => n291, A2 => n290, ZN => O(59));
   U136 : AOI22_X1 port map( A1 => A0(59), A2 => n142, B1 => A4(59), B2 => n173
                           , ZN => n291);
   U137 : AOI222_X1 port map( A1 => A1(59), A2 => n167, B1 => A3(59), B2 => 
                           n159, C1 => A2(59), C2 => n151, ZN => n290);
   U138 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => O(60));
   U139 : AOI22_X1 port map( A1 => A0(60), A2 => n142, B1 => A4(60), B2 => n173
                           , ZN => n295);
   U140 : AOI222_X1 port map( A1 => A1(60), A2 => n167, B1 => A3(60), B2 => 
                           n159, C1 => A2(60), C2 => n151, ZN => n294);
   U141 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => O(61));
   U142 : AOI22_X1 port map( A1 => A0(61), A2 => n142, B1 => A4(61), B2 => n173
                           , ZN => n297);
   U143 : AOI222_X1 port map( A1 => A1(61), A2 => n167, B1 => A3(61), B2 => 
                           n159, C1 => A2(61), C2 => n151, ZN => n296);
   U144 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => O(0));
   U145 : AOI22_X1 port map( A1 => A0(0), A2 => n138, B1 => A4(0), B2 => n178, 
                           ZN => n183);
   U146 : AOI222_X1 port map( A1 => A1(0), A2 => n163, B1 => A3(0), B2 => n155,
                           C1 => A2(0), C2 => n147, ZN => n182);
   U147 : NAND2_X1 port map( A1 => n205, A2 => n204, ZN => O(1));
   U148 : AOI22_X1 port map( A1 => A0(1), A2 => n138, B1 => A4(1), B2 => n177, 
                           ZN => n205);
   U149 : AOI222_X1 port map( A1 => A1(1), A2 => n163, B1 => A3(1), B2 => n155,
                           C1 => A2(1), C2 => n147, ZN => n204);
   U150 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => O(2));
   U151 : AOI22_X1 port map( A1 => A0(2), A2 => n139, B1 => A4(2), B2 => n176, 
                           ZN => n227);
   U152 : AOI222_X1 port map( A1 => A1(2), A2 => n164, B1 => A3(2), B2 => n156,
                           C1 => A2(2), C2 => n148, ZN => n226);
   U153 : NAND2_X1 port map( A1 => n249, A2 => n248, ZN => O(3));
   U154 : AOI22_X1 port map( A1 => A0(3), A2 => n140, B1 => A4(3), B2 => n175, 
                           ZN => n249);
   U155 : AOI222_X1 port map( A1 => A1(3), A2 => n165, B1 => A3(3), B2 => n157,
                           C1 => A2(3), C2 => n149, ZN => n248);
   U156 : NAND2_X1 port map( A1 => n271, A2 => n270, ZN => O(4));
   U157 : AOI22_X1 port map( A1 => A0(4), A2 => n141, B1 => A4(4), B2 => n174, 
                           ZN => n271);
   U158 : AOI222_X1 port map( A1 => A1(4), A2 => n166, B1 => A3(4), B2 => n158,
                           C1 => A2(4), C2 => n150, ZN => n270);
   U159 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => O(5));
   U160 : AOI22_X1 port map( A1 => A0(5), A2 => n142, B1 => A4(5), B2 => n173, 
                           ZN => n293);
   U161 : AOI222_X1 port map( A1 => A1(5), A2 => n167, B1 => A3(5), B2 => n159,
                           C1 => A2(5), C2 => n151, ZN => n292);
   U162 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => O(6));
   U163 : AOI22_X1 port map( A1 => A0(6), A2 => n143, B1 => A4(6), B2 => n173, 
                           ZN => n303);
   U164 : AOI222_X1 port map( A1 => A1(6), A2 => n168, B1 => A3(6), B2 => n160,
                           C1 => A2(6), C2 => n152, ZN => n302);
   U165 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => O(7));
   U166 : AOI22_X1 port map( A1 => A0(7), A2 => n143, B1 => A4(7), B2 => n173, 
                           ZN => n305);
   U167 : AOI222_X1 port map( A1 => A1(7), A2 => n168, B1 => A3(7), B2 => n160,
                           C1 => A2(7), C2 => n152, ZN => n304);
   U168 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => O(8));
   U169 : AOI22_X1 port map( A1 => A0(8), A2 => n143, B1 => A4(8), B2 => n173, 
                           ZN => n307);
   U170 : AOI222_X1 port map( A1 => A1(8), A2 => n168, B1 => A3(8), B2 => n160,
                           C1 => A2(8), C2 => n152, ZN => n306);
   U171 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => O(9));
   U172 : AOI22_X1 port map( A1 => A0(9), A2 => n143, B1 => n178, B2 => A4(9), 
                           ZN => n311);
   U173 : AOI222_X1 port map( A1 => A1(9), A2 => n168, B1 => A3(9), B2 => n160,
                           C1 => A2(9), C2 => n152, ZN => n310);
   U174 : NAND2_X1 port map( A1 => n185, A2 => n184, ZN => O(10));
   U175 : AOI22_X1 port map( A1 => A0(10), A2 => n138, B1 => A4(10), B2 => n178
                           , ZN => n185);
   U176 : AOI222_X1 port map( A1 => A1(10), A2 => n163, B1 => A3(10), B2 => 
                           n155, C1 => A2(10), C2 => n147, ZN => n184);
   U177 : NAND2_X1 port map( A1 => n187, A2 => n186, ZN => O(11));
   U178 : AOI22_X1 port map( A1 => A0(11), A2 => n138, B1 => A4(11), B2 => n178
                           , ZN => n187);
   U179 : AOI222_X1 port map( A1 => A1(11), A2 => n163, B1 => A3(11), B2 => 
                           n155, C1 => A2(11), C2 => n147, ZN => n186);
   U180 : NAND2_X1 port map( A1 => n189, A2 => n188, ZN => O(12));
   U181 : AOI22_X1 port map( A1 => A0(12), A2 => n138, B1 => A4(12), B2 => n177
                           , ZN => n189);
   U182 : AOI222_X1 port map( A1 => A1(12), A2 => n163, B1 => A3(12), B2 => 
                           n155, C1 => A2(12), C2 => n147, ZN => n188);
   U183 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => O(13));
   U184 : AOI22_X1 port map( A1 => A0(13), A2 => n138, B1 => A4(13), B2 => n177
                           , ZN => n191);
   U185 : AOI222_X1 port map( A1 => A1(13), A2 => n163, B1 => A3(13), B2 => 
                           n155, C1 => A2(13), C2 => n147, ZN => n190);
   U186 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => O(14));
   U187 : AOI22_X1 port map( A1 => A0(14), A2 => n138, B1 => A4(14), B2 => n177
                           , ZN => n193);
   U188 : AOI222_X1 port map( A1 => A1(14), A2 => n163, B1 => A3(14), B2 => 
                           n155, C1 => A2(14), C2 => n147, ZN => n192);
   U189 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => O(15));
   U190 : AOI22_X1 port map( A1 => A0(15), A2 => n138, B1 => A4(15), B2 => n177
                           , ZN => n195);
   U191 : AOI222_X1 port map( A1 => A1(15), A2 => n163, B1 => A3(15), B2 => 
                           n155, C1 => A2(15), C2 => n147, ZN => n194);
   U192 : NAND2_X1 port map( A1 => n197, A2 => n196, ZN => O(16));
   U193 : AOI22_X1 port map( A1 => A0(16), A2 => n138, B1 => A4(16), B2 => n177
                           , ZN => n197);
   U194 : AOI222_X1 port map( A1 => A1(16), A2 => n163, B1 => A3(16), B2 => 
                           n155, C1 => A2(16), C2 => n147, ZN => n196);
   U195 : NAND2_X1 port map( A1 => n199, A2 => n198, ZN => O(17));
   U196 : AOI22_X1 port map( A1 => A0(17), A2 => n138, B1 => A4(17), B2 => n177
                           , ZN => n199);
   U197 : AOI222_X1 port map( A1 => A1(17), A2 => n163, B1 => A3(17), B2 => 
                           n155, C1 => A2(17), C2 => n147, ZN => n198);
   U198 : NAND2_X1 port map( A1 => n201, A2 => n200, ZN => O(18));
   U199 : AOI22_X1 port map( A1 => A0(18), A2 => n138, B1 => A4(18), B2 => n177
                           , ZN => n201);
   U200 : AOI222_X1 port map( A1 => A1(18), A2 => n163, B1 => A3(18), B2 => 
                           n155, C1 => A2(18), C2 => n147, ZN => n200);
   U201 : NAND2_X1 port map( A1 => n203, A2 => n202, ZN => O(19));
   U202 : AOI22_X1 port map( A1 => A0(19), A2 => n138, B1 => A4(19), B2 => n177
                           , ZN => n203);
   U203 : AOI222_X1 port map( A1 => A1(19), A2 => n163, B1 => A3(19), B2 => 
                           n155, C1 => A2(19), C2 => n147, ZN => n202);
   U204 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => O(20));
   U205 : AOI22_X1 port map( A1 => A0(20), A2 => n139, B1 => A4(20), B2 => n177
                           , ZN => n207);
   U206 : AOI222_X1 port map( A1 => A1(20), A2 => n164, B1 => A3(20), B2 => 
                           n156, C1 => A2(20), C2 => n148, ZN => n206);
   U207 : NAND2_X1 port map( A1 => n209, A2 => n208, ZN => O(21));
   U208 : AOI22_X1 port map( A1 => A0(21), A2 => n139, B1 => A4(21), B2 => n177
                           , ZN => n209);
   U209 : AOI222_X1 port map( A1 => A1(21), A2 => n164, B1 => A3(21), B2 => 
                           n156, C1 => A2(21), C2 => n148, ZN => n208);
   U210 : NAND2_X1 port map( A1 => n211, A2 => n210, ZN => O(22));
   U211 : AOI22_X1 port map( A1 => A0(22), A2 => n139, B1 => A4(22), B2 => n177
                           , ZN => n211);
   U212 : AOI222_X1 port map( A1 => A1(22), A2 => n164, B1 => A3(22), B2 => 
                           n156, C1 => A2(22), C2 => n148, ZN => n210);
   U213 : NAND2_X1 port map( A1 => n213, A2 => n212, ZN => O(23));
   U214 : AOI22_X1 port map( A1 => A0(23), A2 => n139, B1 => A4(23), B2 => n176
                           , ZN => n213);
   U215 : AOI222_X1 port map( A1 => A1(23), A2 => n164, B1 => A3(23), B2 => 
                           n156, C1 => A2(23), C2 => n148, ZN => n212);
   U216 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => O(24));
   U217 : AOI22_X1 port map( A1 => A0(24), A2 => n139, B1 => A4(24), B2 => n176
                           , ZN => n215);
   U218 : AOI222_X1 port map( A1 => A1(24), A2 => n164, B1 => A3(24), B2 => 
                           n156, C1 => A2(24), C2 => n148, ZN => n214);
   U219 : NAND2_X1 port map( A1 => n217, A2 => n216, ZN => O(25));
   U220 : AOI22_X1 port map( A1 => A0(25), A2 => n139, B1 => A4(25), B2 => n176
                           , ZN => n217);
   U221 : AOI222_X1 port map( A1 => A1(25), A2 => n164, B1 => A3(25), B2 => 
                           n156, C1 => A2(25), C2 => n148, ZN => n216);
   U222 : NAND2_X1 port map( A1 => n219, A2 => n218, ZN => O(26));
   U223 : AOI22_X1 port map( A1 => A0(26), A2 => n139, B1 => A4(26), B2 => n176
                           , ZN => n219);
   U224 : AOI222_X1 port map( A1 => A1(26), A2 => n164, B1 => A3(26), B2 => 
                           n156, C1 => A2(26), C2 => n148, ZN => n218);
   U225 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => O(27));
   U226 : AOI22_X1 port map( A1 => A0(27), A2 => n139, B1 => A4(27), B2 => n176
                           , ZN => n221);
   U227 : AOI222_X1 port map( A1 => A1(27), A2 => n164, B1 => A3(27), B2 => 
                           n156, C1 => A2(27), C2 => n148, ZN => n220);
   U228 : NAND2_X1 port map( A1 => n223, A2 => n222, ZN => O(28));
   U229 : AOI22_X1 port map( A1 => A0(28), A2 => n139, B1 => A4(28), B2 => n176
                           , ZN => n223);
   U230 : AOI222_X1 port map( A1 => A1(28), A2 => n164, B1 => A3(28), B2 => 
                           n156, C1 => A2(28), C2 => n148, ZN => n222);
   U231 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => O(29));
   U232 : AOI22_X1 port map( A1 => A0(29), A2 => n139, B1 => A4(29), B2 => n176
                           , ZN => n225);
   U233 : AOI222_X1 port map( A1 => A1(29), A2 => n164, B1 => A3(29), B2 => 
                           n156, C1 => A2(29), C2 => n148, ZN => n224);
   U234 : AOI222_X1 port map( A1 => A1(39), A2 => n165, B1 => A3(39), B2 => 
                           n157, C1 => A2(39), C2 => n149, ZN => n246);
   U235 : AOI222_X1 port map( A1 => A1(32), A2 => n165, B1 => A3(32), B2 => 
                           n157, C1 => A2(32), C2 => n149, ZN => n232);
   U236 : AOI22_X1 port map( A1 => A0(34), A2 => n140, B1 => A4(34), B2 => n175
                           , ZN => n237);
   U237 : AOI222_X1 port map( A1 => A1(34), A2 => n165, B1 => A3(34), B2 => 
                           n157, C1 => A2(34), C2 => n149, ZN => n236);
   U238 : AOI222_X1 port map( A1 => A1(37), A2 => n165, B1 => A3(37), B2 => 
                           n157, C1 => A2(37), C2 => n149, ZN => n242);
   U239 : AOI222_X1 port map( A1 => A1(33), A2 => n165, B1 => A3(33), B2 => 
                           n157, C1 => A2(33), C2 => n149, ZN => n234);
   U240 : AOI222_X1 port map( A1 => A1(35), A2 => n165, B1 => A3(35), B2 => 
                           n157, C1 => A2(35), C2 => n149, ZN => n238);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_15 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_15;

architecture SYN_BEHAVIORAL of BE_BLOCK_15 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n12, n13 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n12, A2 => n10, B1 => b(2), B2 => n5, ZN => 
                           sel(1));
   U4 : AND2_X1 port map( A1 => n6, A2 => b(2), ZN => n4);
   U5 : AND2_X1 port map( A1 => n12, A2 => n4, ZN => sel(2));
   U6 : AOI21_X1 port map( B1 => n9, B2 => n8, A => b(2), ZN => sel(0));
   U7 : INV_X1 port map( A => b(2), ZN => n10);
   U8 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n5);
   U9 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n6);
   U10 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U11 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n8);
   U12 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n13, ZN => n9);
   U13 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n13);
   U14 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_14 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_14;

architecture SYN_BEHAVIORAL of BE_BLOCK_14 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : INV_X1 port map( A => b(2), ZN => n7);
   U4 : AND3_X1 port map( A1 => b(2), A2 => n4, A3 => n6, ZN => sel(2));
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n4);
   U6 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n5);
   U7 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n4, ZN => n6);
   U8 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n10);
   U9 : AOI21_X1 port map( B1 => n9, B2 => n5, A => b(2), ZN => sel(0));
   U10 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n10, ZN => n9);
   U11 : OAI22_X1 port map( A1 => n7, A2 => n6, B1 => b(2), B2 => n5, ZN => 
                           sel(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_13 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_13;

architecture SYN_BEHAVIORAL of BE_BLOCK_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U4 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U6 : INV_X1 port map( A => b(2), ZN => n4);
   U7 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));
   U8 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_12 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_12;

architecture SYN_BEHAVIORAL of BE_BLOCK_12 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_11 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_11;

architecture SYN_BEHAVIORAL of BE_BLOCK_11 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_10 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_10;

architecture SYN_BEHAVIORAL of BE_BLOCK_10 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_9 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_9;

architecture SYN_BEHAVIORAL of BE_BLOCK_9 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_8 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_8;

architecture SYN_BEHAVIORAL of BE_BLOCK_8 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_7 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_7;

architecture SYN_BEHAVIORAL of BE_BLOCK_7 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_6 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_6;

architecture SYN_BEHAVIORAL of BE_BLOCK_6 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_5 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_5;

architecture SYN_BEHAVIORAL of BE_BLOCK_5 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_4 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_4;

architecture SYN_BEHAVIORAL of BE_BLOCK_4 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_3 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_3;

architecture SYN_BEHAVIORAL of BE_BLOCK_3 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_2 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_2;

architecture SYN_BEHAVIORAL of BE_BLOCK_2 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_1 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_1;

architecture SYN_BEHAVIORAL of BE_BLOCK_1 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => n6, B2 => n7, A => b(2), ZN => sel(0));
   U4 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n7);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => b(2), B2 => n7, ZN => 
                           sel(1));
   U7 : INV_X1 port map( A => b(2), ZN => n4);
   U8 : AND3_X1 port map( A1 => b(2), A2 => n7, A3 => n6, ZN => sel(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BOOTHMUL_DW01_sub_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end BOOTHMUL_DW01_sub_0;

architecture SYN_rpl of BOOTHMUL_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_32_port, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n33, DIFF_9_port, DIFF_12_port, DIFF_13_port, DIFF_15_port, 
      n100, n101, DIFF_6_port, DIFF_31_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, 
      DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, 
      DIFF_29_port, DIFF_30_port, DIFF_7_port, DIFF_5_port, n120, DIFF_4_port, 
      DIFF_11_port, DIFF_8_port, DIFF_10_port, DIFF_14_port, DIFF_16_port, 
      DIFF_3_port, n128, DIFF_1_port, n130, DIFF_2_port, n132, n133, n134, n135
      , n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161 : std_logic;

begin
   DIFF <= ( DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, 
      DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, 
      DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, 
      DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, 
      DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, 
      DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, 
      DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : AND2_X1 port map( A1 => n135, A2 => n130, ZN => n6);
   U2 : XOR2_X1 port map( A => n139, B => n9, Z => DIFF_9_port);
   U3 : XOR2_X1 port map( A => n142, B => n12, Z => DIFF_12_port);
   U4 : XOR2_X1 port map( A => n143, B => n13, Z => DIFF_13_port);
   U5 : XOR2_X1 port map( A => n145, B => n15, Z => DIFF_15_port);
   U6 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n100);
   U7 : AND2_X1 port map( A1 => n100, A2 => n101, ZN => n4);
   U8 : AND2_X1 port map( A1 => n133, A2 => n132, ZN => n101);
   U9 : XOR2_X1 port map( A => n136, B => n6, Z => DIFF_6_port);
   U10 : XNOR2_X1 port map( A => n3, B => B(3), ZN => DIFF_3_port);
   U11 : XOR2_X1 port map( A => n161, B => n31, Z => DIFF_31_port);
   U12 : XOR2_X1 port map( A => n147, B => n17, Z => DIFF_17_port);
   U13 : XOR2_X1 port map( A => n148, B => n18, Z => DIFF_18_port);
   U14 : XOR2_X1 port map( A => n149, B => n19, Z => DIFF_19_port);
   U15 : XOR2_X1 port map( A => n150, B => n20, Z => DIFF_20_port);
   U16 : XOR2_X1 port map( A => n151, B => n21, Z => DIFF_21_port);
   U17 : XOR2_X1 port map( A => n152, B => n22, Z => DIFF_22_port);
   U18 : XOR2_X1 port map( A => n153, B => n23, Z => DIFF_23_port);
   U19 : XOR2_X1 port map( A => n154, B => n24, Z => DIFF_24_port);
   U20 : XOR2_X1 port map( A => n155, B => n25, Z => DIFF_25_port);
   U21 : XOR2_X1 port map( A => n156, B => n26, Z => DIFF_26_port);
   U22 : XOR2_X1 port map( A => n157, B => n27, Z => DIFF_27_port);
   U23 : XOR2_X1 port map( A => n158, B => n28, Z => DIFF_28_port);
   U24 : XOR2_X1 port map( A => n159, B => n29, Z => DIFF_29_port);
   U25 : XOR2_X1 port map( A => n160, B => n30, Z => DIFF_30_port);
   U26 : XNOR2_X1 port map( A => n161, B => n33, ZN => DIFF_32_port);
   U27 : NAND2_X1 port map( A1 => n161, A2 => n31, ZN => n33);
   U28 : XOR2_X1 port map( A => n137, B => n7, Z => DIFF_7_port);
   U29 : AND2_X1 port map( A1 => n136, A2 => n6, ZN => n7);
   U30 : XNOR2_X1 port map( A => n120, B => n135, ZN => DIFF_5_port);
   U31 : NAND2_X1 port map( A1 => n134, A2 => n4, ZN => n120);
   U32 : XOR2_X1 port map( A => n134, B => n4, Z => DIFF_4_port);
   U33 : XOR2_X1 port map( A => n141, B => n11, Z => DIFF_11_port);
   U34 : XOR2_X1 port map( A => n138, B => n8, Z => DIFF_8_port);
   U35 : AND2_X1 port map( A1 => n137, A2 => n7, ZN => n8);
   U36 : AND2_X1 port map( A1 => n148, A2 => n18, ZN => n19);
   U37 : AND2_X1 port map( A1 => n147, A2 => n17, ZN => n18);
   U38 : AND2_X1 port map( A1 => n146, A2 => n16, ZN => n17);
   U39 : AND2_X1 port map( A1 => n145, A2 => n15, ZN => n16);
   U40 : AND2_X1 port map( A1 => n144, A2 => n14, ZN => n15);
   U41 : AND2_X1 port map( A1 => n143, A2 => n13, ZN => n14);
   U42 : AND2_X1 port map( A1 => n142, A2 => n12, ZN => n13);
   U43 : AND2_X1 port map( A1 => n141, A2 => n11, ZN => n12);
   U44 : AND2_X1 port map( A1 => n149, A2 => n19, ZN => n20);
   U45 : AND2_X1 port map( A1 => n138, A2 => n8, ZN => n9);
   U46 : AND2_X1 port map( A1 => n150, A2 => n20, ZN => n21);
   U47 : XOR2_X1 port map( A => n140, B => n10, Z => DIFF_10_port);
   U48 : AND2_X1 port map( A1 => n139, A2 => n9, ZN => n10);
   U49 : XOR2_X1 port map( A => n144, B => n14, Z => DIFF_14_port);
   U50 : AND2_X1 port map( A1 => n151, A2 => n21, ZN => n22);
   U51 : AND2_X1 port map( A1 => n140, A2 => n10, ZN => n11);
   U52 : AND2_X1 port map( A1 => n160, A2 => n30, ZN => n31);
   U53 : AND2_X1 port map( A1 => n159, A2 => n29, ZN => n30);
   U54 : AND2_X1 port map( A1 => n158, A2 => n28, ZN => n29);
   U55 : AND2_X1 port map( A1 => n157, A2 => n27, ZN => n28);
   U56 : AND2_X1 port map( A1 => n156, A2 => n26, ZN => n27);
   U57 : AND2_X1 port map( A1 => n155, A2 => n25, ZN => n26);
   U58 : AND2_X1 port map( A1 => n154, A2 => n24, ZN => n25);
   U59 : AND2_X1 port map( A1 => n153, A2 => n23, ZN => n24);
   U60 : AND2_X1 port map( A1 => n152, A2 => n22, ZN => n23);
   U61 : XOR2_X1 port map( A => n146, B => n16, Z => DIFF_16_port);
   U62 : INV_X1 port map( A => B(32), ZN => n161);
   U63 : INV_X1 port map( A => B(11), ZN => n141);
   U64 : INV_X1 port map( A => B(12), ZN => n142);
   U65 : INV_X1 port map( A => B(13), ZN => n143);
   U66 : INV_X1 port map( A => B(14), ZN => n144);
   U67 : INV_X1 port map( A => B(15), ZN => n145);
   U68 : INV_X1 port map( A => B(16), ZN => n146);
   U69 : INV_X1 port map( A => B(17), ZN => n147);
   U70 : INV_X1 port map( A => B(18), ZN => n148);
   U71 : INV_X1 port map( A => B(19), ZN => n149);
   U72 : INV_X1 port map( A => B(20), ZN => n150);
   U73 : INV_X1 port map( A => B(21), ZN => n151);
   U74 : INV_X1 port map( A => B(22), ZN => n152);
   U75 : INV_X1 port map( A => B(23), ZN => n153);
   U76 : INV_X1 port map( A => B(24), ZN => n154);
   U77 : INV_X1 port map( A => B(25), ZN => n155);
   U78 : INV_X1 port map( A => B(26), ZN => n156);
   U79 : INV_X1 port map( A => B(27), ZN => n157);
   U80 : INV_X1 port map( A => B(28), ZN => n158);
   U81 : INV_X1 port map( A => B(29), ZN => n159);
   U82 : INV_X1 port map( A => B(30), ZN => n160);
   U83 : AND2_X1 port map( A1 => n2, A2 => n132, ZN => n3);
   U84 : NOR2_X1 port map( A1 => B(1), A2 => B(0), ZN => n128);
   U85 : NOR2_X1 port map( A1 => B(1), A2 => B(0), ZN => n2);
   U86 : INV_X1 port map( A => B(10), ZN => n140);
   U87 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U88 : AND2_X1 port map( A1 => n134, A2 => n4, ZN => n130);
   U89 : INV_X1 port map( A => B(9), ZN => n139);
   U90 : INV_X1 port map( A => B(7), ZN => n137);
   U91 : XNOR2_X1 port map( A => B(2), B => n128, ZN => DIFF_2_port);
   U92 : INV_X1 port map( A => B(8), ZN => n138);
   U93 : INV_X1 port map( A => B(2), ZN => n132);
   U94 : INV_X1 port map( A => B(6), ZN => n136);
   U95 : INV_X1 port map( A => B(5), ZN => n135);
   U96 : INV_X1 port map( A => B(4), ZN => n134);
   U97 : INV_X1 port map( A => B(3), ZN => n133);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NBIT64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_0;

architecture SYN_STRUCTURAL of RCA_NBIT64_0 is

   component FA_897
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_898
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_899
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_900
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_901
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_902
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_903
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_904
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_905
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_906
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_907
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_908
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_909
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_910
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_911
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_912
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_913
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_914
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_915
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_916
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_917
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_918
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_919
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_959 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_958 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_957 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_956 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_955 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_954 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_953 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_952 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_951 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_950 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_949 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_948 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_947 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_946 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_945 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_944 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_943 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_942 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_941 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_940 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_939 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_938 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_937 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_936 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_935 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_934 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_933 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_932 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_931 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_930 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_929 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_928 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_927 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_926 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_925 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_924 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_923 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_922 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_921 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_920 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_919 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_918 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_917 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_916 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_915 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_914 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_913 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_912 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_911 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_910 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_909 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_908 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_907 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_906 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_905 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_904 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_903 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_902 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_901 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_900 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_899 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_898 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_897 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX_5TO1_NBIT64_0 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX_5TO1_NBIT64_0;

architecture SYN_BEHAVIORAL of MUX_5TO1_NBIT64_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, net127215, net127213, net127211, net127203, net127217, 
      net127229, net127227, net127225, net127219, net129570, net129567, 
      net129583, net129581, net129580, net129752, net129805, net129799, 
      net129797, net129793, net129791, net129807, net129941, net129937, 
      net129955, net129947, net129945, net131633, net136967, net137140, 
      net137139, net137138, net153432, net137097, net137096, net136985, 
      net136172, n89, n88, n5, net137098, n6, n136, n137, n138, n139, n140 : 
      std_logic;

begin
   
   U1 : BUF_X4 port map( A => net129580, Z => net129583);
   U2 : CLKBUF_X1 port map( A => net127203, Z => net129941);
   U3 : BUF_X4 port map( A => net129941, Z => net129937);
   U4 : BUF_X2 port map( A => net129955, Z => net129945);
   U5 : BUF_X2 port map( A => net129567, Z => net129570);
   U6 : CLKBUF_X1 port map( A => net129807, Z => net129805);
   U7 : BUF_X2 port map( A => net129805, Z => net129791);
   U8 : CLKBUF_X1 port map( A => net129791, Z => net129797);
   U9 : CLKBUF_X1 port map( A => net131633, Z => net127229);
   U10 : CLKBUF_X1 port map( A => net131633, Z => net127227);
   U11 : CLKBUF_X1 port map( A => net131633, Z => net127225);
   U12 : BUF_X1 port map( A => net127215, Z => net127203);
   U13 : AND2_X1 port map( A1 => A2(2), A2 => n6, ZN => net137098);
   U14 : NOR3_X1 port map( A1 => net137097, A2 => net137096, A3 => net137098, 
                           ZN => n89);
   U15 : AND2_X1 port map( A1 => sel(1), A2 => n136, ZN => n6);
   U16 : CLKBUF_X1 port map( A => n6, Z => net127217);
   U17 : AND2_X1 port map( A1 => A2(3), A2 => n6, ZN => net137140);
   U18 : INV_X1 port map( A => sel(0), ZN => n136);
   U19 : NOR2_X1 port map( A1 => sel(1), A2 => n136, ZN => net153432);
   U20 : AND2_X1 port map( A1 => net136172, A2 => sel(1), ZN => n5);
   U21 : CLKBUF_X1 port map( A => sel(1), Z => net136967);
   U22 : BUF_X1 port map( A => sel(0), Z => net136172);
   U23 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => O(2));
   U24 : AND2_X1 port map( A1 => A1(2), A2 => net153432, ZN => net137096);
   U25 : AND2_X1 port map( A1 => A3(2), A2 => n5, ZN => net137097);
   U26 : AOI22_X1 port map( A1 => A0(2), A2 => net131633, B1 => A4(2), B2 => 
                           n137, ZN => n88);
   U27 : CLKBUF_X1 port map( A => sel(2), Z => n137);
   U28 : AOI22_X1 port map( A1 => A0(9), A2 => net127229, B1 => n137, B2 => 
                           A4(9), ZN => n2);
   U29 : AOI22_X1 port map( A1 => A0(3), A2 => net131633, B1 => A4(3), B2 => 
                           n137, ZN => n66);
   U30 : AOI22_X1 port map( A1 => A0(5), A2 => net127227, B1 => A4(5), B2 => 
                           n137, ZN => n22);
   U31 : BUF_X1 port map( A => net127225, Z => net127219);
   U32 : BUF_X2 port map( A => net153432, Z => net129580);
   U33 : AND2_X1 port map( A1 => A1(3), A2 => net153432, ZN => net137138);
   U34 : CLKBUF_X1 port map( A => n5, Z => net129567);
   U35 : AND2_X1 port map( A1 => A3(3), A2 => n5, ZN => net137139);
   U36 : CLKBUF_X1 port map( A => net136172, Z => net136985);
   U37 : CLKBUF_X1 port map( A => sel(2), Z => net129807);
   U38 : NOR3_X1 port map( A1 => net136967, A2 => net129799, A3 => net136985, 
                           ZN => net131633);
   U39 : NOR3_X1 port map( A1 => net137138, A2 => net137139, A3 => net137140, 
                           ZN => n67);
   U40 : BUF_X2 port map( A => net129945, Z => net129947);
   U41 : BUF_X1 port map( A => net127217, Z => net127215);
   U42 : BUF_X1 port map( A => net129805, Z => net129793);
   U43 : BUF_X1 port map( A => net129807, Z => net129799);
   U44 : AOI22_X1 port map( A1 => A0(7), A2 => net127229, B1 => A4(7), B2 => 
                           net129793, ZN => n10);
   U45 : AOI22_X1 port map( A1 => A0(11), A2 => net127219, B1 => A4(11), B2 => 
                           net129791, ZN => n128);
   U46 : AOI222_X1 port map( A1 => A1(11), A2 => net129581, B1 => A3(11), B2 =>
                           net129570, C1 => A2(11), C2 => net127211, ZN => n129
                           );
   U47 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => O(8));
   U48 : AOI22_X1 port map( A1 => A0(8), A2 => net127229, B1 => A4(8), B2 => 
                           net129793, ZN => n8);
   U49 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => O(19));
   U50 : AOI22_X1 port map( A1 => A0(19), A2 => net127219, B1 => A4(19), B2 => 
                           net129791, ZN => n112);
   U51 : AOI222_X1 port map( A1 => A1(19), A2 => net129583, B1 => A3(19), B2 =>
                           net129947, C1 => A2(19), C2 => net129937, ZN => n113
                           );
   U52 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => O(18));
   U53 : AOI22_X1 port map( A1 => A0(18), A2 => net127219, B1 => A4(18), B2 => 
                           net129791, ZN => n114);
   U54 : AOI22_X1 port map( A1 => A0(12), A2 => net127219, B1 => A4(12), B2 => 
                           net129791, ZN => n126);
   U55 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => O(20));
   U56 : AOI22_X1 port map( A1 => A0(20), A2 => net127229, B1 => A4(20), B2 => 
                           net129791, ZN => n108);
   U57 : AOI222_X1 port map( A1 => A1(20), A2 => net129752, B1 => A3(20), B2 =>
                           net129947, C1 => A2(20), C2 => net129937, ZN => n109
                           );
   U58 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => O(17));
   U59 : AOI22_X1 port map( A1 => A0(17), A2 => net127219, B1 => A4(17), B2 => 
                           net129791, ZN => n116);
   U60 : AOI22_X1 port map( A1 => A0(13), A2 => net127219, B1 => A4(13), B2 => 
                           net129793, ZN => n124);
   U61 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => O(21));
   U62 : AOI22_X1 port map( A1 => A0(21), A2 => net127227, B1 => A4(21), B2 => 
                           net129791, ZN => n106);
   U63 : AOI222_X1 port map( A1 => A1(21), A2 => net129583, B1 => A3(21), B2 =>
                           net129947, C1 => A2(21), C2 => net129937, ZN => n107
                           );
   U64 : AOI22_X1 port map( A1 => A0(16), A2 => net127219, B1 => A4(16), B2 => 
                           net129791, ZN => n118);
   U65 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => O(10));
   U66 : AOI22_X1 port map( A1 => A0(10), A2 => net127219, B1 => A4(10), B2 => 
                           net129791, ZN => n130);
   U67 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => O(15));
   U68 : AOI22_X1 port map( A1 => A0(15), A2 => net127219, B1 => A4(15), B2 => 
                           net129791, ZN => n120);
   U69 : AOI22_X1 port map( A1 => A0(14), A2 => net127219, B1 => A4(14), B2 => 
                           net129791, ZN => n122);
   U70 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => O(22));
   U71 : AOI22_X1 port map( A1 => A0(22), A2 => net127227, B1 => A4(22), B2 => 
                           net129791, ZN => n104);
   U72 : AOI222_X1 port map( A1 => A1(22), A2 => net129580, B1 => A3(22), B2 =>
                           net129947, C1 => A2(22), C2 => net129937, ZN => n105
                           );
   U73 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => O(32));
   U74 : AOI22_X1 port map( A1 => A0(32), A2 => net127227, B1 => A4(32), B2 => 
                           net129797, ZN => n82);
   U75 : AOI222_X1 port map( A1 => A1(32), A2 => net129752, B1 => A3(32), B2 =>
                           net129947, C1 => A2(32), C2 => net129937, ZN => n83)
                           ;
   U76 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => O(23));
   U77 : AOI22_X1 port map( A1 => A0(23), A2 => net127227, B1 => A4(23), B2 => 
                           net129793, ZN => n102);
   U78 : AOI222_X1 port map( A1 => A1(23), A2 => net129581, B1 => A3(23), B2 =>
                           net129947, C1 => A2(23), C2 => net129937, ZN => n103
                           );
   U79 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => O(24));
   U80 : AOI22_X1 port map( A1 => A0(24), A2 => net127227, B1 => A4(24), B2 => 
                           net129793, ZN => n100);
   U81 : AOI222_X1 port map( A1 => A1(24), A2 => net129752, B1 => A3(24), B2 =>
                           net129947, C1 => A2(24), C2 => net129937, ZN => n101
                           );
   U82 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => O(33));
   U83 : AOI22_X1 port map( A1 => A0(33), A2 => net127225, B1 => A4(33), B2 => 
                           net129799, ZN => n80);
   U84 : AOI222_X1 port map( A1 => A1(33), A2 => net129583, B1 => A3(33), B2 =>
                           net129947, C1 => A2(33), C2 => net129937, ZN => n81)
                           ;
   U85 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => O(25));
   U86 : AOI22_X1 port map( A1 => A0(25), A2 => net127227, B1 => A4(25), B2 => 
                           net129793, ZN => n98);
   U87 : AOI222_X1 port map( A1 => A1(25), A2 => net129583, B1 => A3(25), B2 =>
                           net129947, C1 => A2(25), C2 => net129937, ZN => n99)
                           ;
   U88 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => O(26));
   U89 : AOI22_X1 port map( A1 => A0(26), A2 => net127227, B1 => A4(26), B2 => 
                           net129791, ZN => n96);
   U90 : AOI222_X1 port map( A1 => A1(26), A2 => net129752, B1 => A3(26), B2 =>
                           net129947, C1 => A2(26), C2 => net129937, ZN => n97)
                           ;
   U91 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => O(34));
   U92 : AOI22_X1 port map( A1 => A0(34), A2 => net127225, B1 => A4(34), B2 => 
                           net129799, ZN => n78);
   U93 : AOI222_X1 port map( A1 => A1(34), A2 => net129580, B1 => A3(34), B2 =>
                           net129947, C1 => A2(34), C2 => net129937, ZN => n79)
                           ;
   U94 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => O(27));
   U95 : AOI22_X1 port map( A1 => A0(27), A2 => net127229, B1 => A4(27), B2 => 
                           net129797, ZN => n94);
   U96 : AOI222_X1 port map( A1 => A1(27), A2 => net129583, B1 => A3(27), B2 =>
                           net129947, C1 => A2(27), C2 => net129937, ZN => n95)
                           ;
   U97 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => O(28));
   U98 : AOI22_X1 port map( A1 => A0(28), A2 => net127227, B1 => A4(28), B2 => 
                           net129799, ZN => n92);
   U99 : AOI222_X1 port map( A1 => A1(28), A2 => net129580, B1 => A3(28), B2 =>
                           net129947, C1 => A2(28), C2 => net129937, ZN => n93)
                           ;
   U100 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => O(29));
   U101 : AOI22_X1 port map( A1 => A0(29), A2 => net127229, B1 => A4(29), B2 =>
                           net129799, ZN => n90);
   U102 : AOI222_X1 port map( A1 => A1(29), A2 => net129581, B1 => A3(29), B2 
                           => net129947, C1 => A2(29), C2 => net129937, ZN => 
                           n91);
   U103 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => O(35));
   U104 : AOI22_X1 port map( A1 => A0(35), A2 => net127219, B1 => A4(35), B2 =>
                           net129799, ZN => n76);
   U105 : AOI222_X1 port map( A1 => A1(35), A2 => net129581, B1 => A3(35), B2 
                           => net129947, C1 => A2(35), C2 => net129937, ZN => 
                           n77);
   U106 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => O(30));
   U107 : AOI22_X1 port map( A1 => A0(30), A2 => net127229, B1 => A4(30), B2 =>
                           net129799, ZN => n86);
   U108 : AOI222_X1 port map( A1 => A1(30), A2 => net129752, B1 => A3(30), B2 
                           => net129947, C1 => A2(30), C2 => net129937, ZN => 
                           n87);
   U109 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => O(31));
   U110 : AOI22_X1 port map( A1 => A0(31), A2 => net127229, B1 => A4(31), B2 =>
                           net129799, ZN => n84);
   U111 : AOI222_X1 port map( A1 => A1(31), A2 => net129583, B1 => A3(31), B2 
                           => net129947, C1 => A2(31), C2 => net129937, ZN => 
                           n85);
   U112 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => O(36));
   U113 : AOI22_X1 port map( A1 => A0(36), A2 => net127227, B1 => A4(36), B2 =>
                           net129799, ZN => n74);
   U114 : AOI222_X1 port map( A1 => A1(36), A2 => net129752, B1 => A3(36), B2 
                           => net129947, C1 => A2(36), C2 => net129937, ZN => 
                           n75);
   U115 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => O(37));
   U116 : AOI22_X1 port map( A1 => A0(37), A2 => net127229, B1 => A4(37), B2 =>
                           net129799, ZN => n72);
   U117 : AOI222_X1 port map( A1 => A1(37), A2 => net129583, B1 => A3(37), B2 
                           => net129947, C1 => A2(37), C2 => net129937, ZN => 
                           n73);
   U118 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => O(38));
   U119 : AOI22_X1 port map( A1 => A0(38), A2 => net127229, B1 => A4(38), B2 =>
                           net129797, ZN => n70);
   U120 : AOI222_X1 port map( A1 => A1(38), A2 => net129752, B1 => A3(38), B2 
                           => net129947, C1 => A2(38), C2 => net129937, ZN => 
                           n71);
   U121 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => O(39));
   U122 : AOI22_X1 port map( A1 => A0(39), A2 => net127227, B1 => A4(39), B2 =>
                           net129799, ZN => n68);
   U123 : AOI222_X1 port map( A1 => A1(39), A2 => net129583, B1 => A3(39), B2 
                           => net129947, C1 => A2(39), C2 => net129937, ZN => 
                           n69);
   U124 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => O(40));
   U125 : AOI22_X1 port map( A1 => A0(40), A2 => net127229, B1 => A4(40), B2 =>
                           net129797, ZN => n64);
   U126 : AOI222_X1 port map( A1 => A1(40), A2 => net129580, B1 => A3(40), B2 
                           => net129947, C1 => A2(40), C2 => net129937, ZN => 
                           n65);
   U127 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => O(41));
   U128 : AOI22_X1 port map( A1 => A0(41), A2 => net127227, B1 => A4(41), B2 =>
                           net129797, ZN => n62);
   U129 : AOI222_X1 port map( A1 => A1(41), A2 => net129581, B1 => A3(41), B2 
                           => net129947, C1 => A2(41), C2 => net129937, ZN => 
                           n63);
   U130 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => O(42));
   U131 : AOI22_X1 port map( A1 => A0(42), A2 => net127225, B1 => A4(42), B2 =>
                           net129797, ZN => n60);
   U132 : AOI222_X1 port map( A1 => A1(42), A2 => net129752, B1 => A3(42), B2 
                           => net129947, C1 => A2(42), C2 => net129937, ZN => 
                           n61);
   U133 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => O(43));
   U134 : AOI22_X1 port map( A1 => A0(43), A2 => net127225, B1 => A4(43), B2 =>
                           net129797, ZN => n58);
   U135 : AOI222_X1 port map( A1 => A1(43), A2 => net129583, B1 => A3(43), B2 
                           => net129947, C1 => A2(43), C2 => net129937, ZN => 
                           n59);
   U136 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => O(44));
   U137 : AOI22_X1 port map( A1 => A0(44), A2 => net127225, B1 => A4(44), B2 =>
                           net129797, ZN => n56);
   U138 : AOI222_X1 port map( A1 => A1(44), A2 => net129752, B1 => A3(44), B2 
                           => net129947, C1 => A2(44), C2 => net129937, ZN => 
                           n57);
   U139 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => O(45));
   U140 : AOI22_X1 port map( A1 => A0(45), A2 => net127225, B1 => A4(45), B2 =>
                           net129797, ZN => n54);
   U141 : AOI222_X1 port map( A1 => A1(45), A2 => net129583, B1 => A3(45), B2 
                           => net129947, C1 => A2(45), C2 => net129937, ZN => 
                           n55);
   U142 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => O(46));
   U143 : AOI22_X1 port map( A1 => A0(46), A2 => net127225, B1 => A4(46), B2 =>
                           net129797, ZN => n52);
   U144 : AOI222_X1 port map( A1 => A1(46), A2 => net129580, B1 => A3(46), B2 
                           => net129947, C1 => A2(46), C2 => net129937, ZN => 
                           n53);
   U145 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => O(47));
   U146 : AOI22_X1 port map( A1 => A0(47), A2 => net127225, B1 => A4(47), B2 =>
                           net129797, ZN => n50);
   U147 : AOI222_X1 port map( A1 => A1(47), A2 => net129581, B1 => A3(47), B2 
                           => net129947, C1 => A2(47), C2 => net129937, ZN => 
                           n51);
   U148 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => O(48));
   U149 : AOI22_X1 port map( A1 => A0(48), A2 => net127225, B1 => A4(48), B2 =>
                           net129797, ZN => n48);
   U150 : AOI222_X1 port map( A1 => A1(48), A2 => net129752, B1 => A3(48), B2 
                           => net129947, C1 => A2(48), C2 => net129937, ZN => 
                           n49);
   U151 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => O(49));
   U152 : AOI22_X1 port map( A1 => A0(49), A2 => net127225, B1 => A4(49), B2 =>
                           net129797, ZN => n46);
   U153 : AOI222_X1 port map( A1 => A1(49), A2 => net129583, B1 => A3(49), B2 
                           => net129947, C1 => A2(49), C2 => net129937, ZN => 
                           n47);
   U154 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => O(50));
   U155 : AOI22_X1 port map( A1 => A0(50), A2 => net127225, B1 => A4(50), B2 =>
                           net129797, ZN => n42);
   U156 : AOI222_X1 port map( A1 => A1(50), A2 => net129752, B1 => A3(50), B2 
                           => net129947, C1 => A2(50), C2 => net129937, ZN => 
                           n43);
   U157 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => O(51));
   U158 : AOI22_X1 port map( A1 => A0(51), A2 => net127225, B1 => A4(51), B2 =>
                           net129797, ZN => n40);
   U159 : AOI222_X1 port map( A1 => A1(51), A2 => net129583, B1 => A3(51), B2 
                           => net129947, C1 => A2(51), C2 => net129937, ZN => 
                           n41);
   U160 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => O(52));
   U161 : AOI22_X1 port map( A1 => A0(52), A2 => net127225, B1 => A4(52), B2 =>
                           net129797, ZN => n38);
   U162 : AOI222_X1 port map( A1 => A1(52), A2 => net129580, B1 => A3(52), B2 
                           => net129947, C1 => A2(52), C2 => net129937, ZN => 
                           n39);
   U163 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => O(53));
   U164 : AOI22_X1 port map( A1 => A0(53), A2 => net127227, B1 => A4(53), B2 =>
                           net129797, ZN => n36);
   U165 : AOI222_X1 port map( A1 => A1(53), A2 => net129581, B1 => A3(53), B2 
                           => net129947, C1 => A2(53), C2 => net129937, ZN => 
                           n37);
   U166 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => O(54));
   U167 : AOI22_X1 port map( A1 => A0(54), A2 => net127227, B1 => A4(54), B2 =>
                           net129797, ZN => n34);
   U168 : AOI222_X1 port map( A1 => A1(54), A2 => net129752, B1 => A3(54), B2 
                           => net129947, C1 => A2(54), C2 => net129937, ZN => 
                           n35);
   U169 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => O(55));
   U170 : AOI22_X1 port map( A1 => A0(55), A2 => net127227, B1 => A4(55), B2 =>
                           net129797, ZN => n32);
   U171 : AOI222_X1 port map( A1 => A1(55), A2 => net129583, B1 => A3(55), B2 
                           => net129947, C1 => A2(55), C2 => net129937, ZN => 
                           n33);
   U172 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => O(56));
   U173 : AOI22_X1 port map( A1 => A0(56), A2 => net127227, B1 => A4(56), B2 =>
                           net129797, ZN => n30);
   U174 : AOI222_X1 port map( A1 => A1(56), A2 => net129752, B1 => A3(56), B2 
                           => net129947, C1 => A2(56), C2 => net129937, ZN => 
                           n31);
   U175 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => O(57));
   U176 : AOI22_X1 port map( A1 => A0(57), A2 => net127227, B1 => A4(57), B2 =>
                           net129797, ZN => n28);
   U177 : AOI222_X1 port map( A1 => A1(57), A2 => net129583, B1 => A3(57), B2 
                           => net129947, C1 => A2(57), C2 => net129937, ZN => 
                           n29);
   U178 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => O(58));
   U179 : AOI22_X1 port map( A1 => A0(58), A2 => net127227, B1 => A4(58), B2 =>
                           net129797, ZN => n26);
   U180 : AOI222_X1 port map( A1 => A1(58), A2 => net129580, B1 => A3(58), B2 
                           => net129947, C1 => A2(58), C2 => net129937, ZN => 
                           n27);
   U181 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => O(59));
   U182 : AOI22_X1 port map( A1 => A0(59), A2 => net127227, B1 => A4(59), B2 =>
                           net129797, ZN => n24);
   U183 : AOI222_X1 port map( A1 => A1(59), A2 => net129581, B1 => A3(59), B2 
                           => net129947, C1 => A2(59), C2 => net129937, ZN => 
                           n25);
   U184 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => O(60));
   U185 : AOI22_X1 port map( A1 => A0(60), A2 => net127227, B1 => A4(60), B2 =>
                           net129793, ZN => n20);
   U186 : AOI222_X1 port map( A1 => A1(60), A2 => net129752, B1 => A3(60), B2 
                           => net129947, C1 => A2(60), C2 => net129937, ZN => 
                           n21);
   U187 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => O(61));
   U188 : AOI22_X1 port map( A1 => A0(61), A2 => net127227, B1 => A4(61), B2 =>
                           net129793, ZN => n18);
   U189 : AOI222_X1 port map( A1 => A1(61), A2 => net129583, B1 => A3(61), B2 
                           => net129947, C1 => A2(61), C2 => net129937, ZN => 
                           n19);
   U190 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => O(62));
   U191 : AOI22_X1 port map( A1 => A0(62), A2 => net127227, B1 => A4(62), B2 =>
                           net129793, ZN => n16);
   U192 : AOI222_X1 port map( A1 => A1(62), A2 => net129580, B1 => A3(62), B2 
                           => net129947, C1 => A2(62), C2 => net129937, ZN => 
                           n17);
   U193 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => O(63));
   U194 : AOI22_X1 port map( A1 => A0(63), A2 => net127227, B1 => A4(63), B2 =>
                           net129793, ZN => n14);
   U195 : AOI222_X1 port map( A1 => A1(63), A2 => net129581, B1 => A3(63), B2 
                           => net129947, C1 => A2(63), C2 => net129937, ZN => 
                           n15);
   U196 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => O(1));
   U197 : AOI22_X1 port map( A1 => A0(1), A2 => net127219, B1 => A4(1), B2 => 
                           net129793, ZN => n110);
   U198 : AOI222_X1 port map( A1 => A1(1), A2 => net129583, B1 => A3(1), B2 => 
                           net129947, C1 => A2(1), C2 => net129937, ZN => n111)
                           ;
   U199 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => O(0));
   U200 : AOI22_X1 port map( A1 => A0(0), A2 => net127219, B1 => A4(0), B2 => 
                           net129793, ZN => n132);
   U201 : AOI222_X1 port map( A1 => A1(0), A2 => net129752, B1 => A3(0), B2 => 
                           net129947, C1 => A2(0), C2 => net129937, ZN => n133)
                           ;
   U202 : AOI222_X1 port map( A1 => A1(18), A2 => net129752, B1 => A3(18), B2 
                           => net129947, C1 => A2(18), C2 => net129937, ZN => 
                           n115);
   U203 : CLKBUF_X1 port map( A => net129570, Z => net129955);
   U204 : CLKBUF_X1 port map( A => net129583, Z => net129752);
   U205 : AOI222_X1 port map( A1 => A1(17), A2 => net129581, B1 => A3(17), B2 
                           => net129945, C1 => A2(17), C2 => net129941, ZN => 
                           n117);
   U206 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => O(16));
   U207 : AOI222_X1 port map( A1 => A1(16), A2 => net129580, B1 => A3(16), B2 
                           => net129945, C1 => A2(16), C2 => net129941, ZN => 
                           n119);
   U208 : AOI222_X1 port map( A1 => A1(15), A2 => net129583, B1 => A3(15), B2 
                           => net129945, C1 => A2(15), C2 => net127203, ZN => 
                           n121);
   U209 : CLKBUF_X1 port map( A => net127217, Z => net127213);
   U210 : BUF_X1 port map( A => net127213, Z => net127211);
   U211 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => O(14));
   U212 : AOI222_X1 port map( A1 => A1(14), A2 => net129583, B1 => A3(14), B2 
                           => net129945, C1 => A2(14), C2 => net127203, ZN => 
                           n123);
   U213 : AOI222_X1 port map( A1 => A1(4), A2 => net129580, B1 => A3(4), B2 => 
                           net129567, C1 => A2(4), C2 => net127217, ZN => n45);
   U214 : BUF_X1 port map( A => net129580, Z => net129581);
   U215 : NAND2_X1 port map( A1 => A1(6), A2 => net129583, ZN => n138);
   U216 : NAND2_X1 port map( A1 => A3(6), A2 => net129570, ZN => n139);
   U217 : NAND2_X1 port map( A1 => A2(6), A2 => net127215, ZN => n140);
   U218 : AND3_X1 port map( A1 => n138, A2 => n139, A3 => n140, ZN => n13);
   U219 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => O(13));
   U220 : AOI222_X1 port map( A1 => A1(13), A2 => net129583, B1 => A3(13), B2 
                           => net129945, C1 => A2(13), C2 => net127203, ZN => 
                           n125);
   U221 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => O(12));
   U222 : AOI222_X1 port map( A1 => A1(12), A2 => net129752, B1 => A3(12), B2 
                           => net129955, C1 => A2(12), C2 => net127203, ZN => 
                           n127);
   U223 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => O(11));
   U224 : AOI222_X1 port map( A1 => A1(10), A2 => net129580, B1 => A3(10), B2 
                           => net129570, C1 => A2(10), C2 => net127211, ZN => 
                           n131);
   U225 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => O(9));
   U226 : AOI222_X1 port map( A1 => A1(9), A2 => net129583, B1 => A3(9), B2 => 
                           net129570, C1 => A2(9), C2 => net127211, ZN => n3);
   U227 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => O(6));
   U228 : AOI22_X1 port map( A1 => A0(6), A2 => net127229, B1 => A4(6), B2 => 
                           net129799, ZN => n12);
   U229 : AOI222_X1 port map( A1 => A1(8), A2 => net129583, B1 => A3(8), B2 => 
                           net129570, C1 => A2(8), C2 => net127215, ZN => n9);
   U230 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => O(7));
   U231 : AOI222_X1 port map( A1 => A1(7), A2 => net129583, B1 => A3(7), B2 => 
                           net129570, C1 => A2(7), C2 => net127213, ZN => n11);
   U232 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => O(5));
   U233 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => O(3));
   U234 : AOI222_X1 port map( A1 => A1(5), A2 => net129581, B1 => A3(5), B2 => 
                           net129570, C1 => A2(5), C2 => net127215, ZN => n23);
   U235 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => O(4));
   U236 : AOI22_X1 port map( A1 => A0(4), A2 => net127225, B1 => A4(4), B2 => 
                           net129799, ZN => n44);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BE_BLOCK_0 is

   port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2 
         downto 0));

end BE_BLOCK_0;

architecture SYN_BEHAVIORAL of BE_BLOCK_0 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net153327, net136198, net125371, n2, n4, n5 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n4);
   U4 : OAI22_X1 port map( A1 => n4, A2 => net125371, B1 => b(2), B2 => n2, ZN 
                           => sel(1));
   U5 : NOR2_X1 port map( A1 => b(1), A2 => b(0), ZN => net153327);
   U6 : BUF_X1 port map( A => b(1), Z => n5);
   U7 : NAND2_X1 port map( A1 => n5, A2 => b(0), ZN => n2);
   U8 : XNOR2_X1 port map( A => n5, B => b(0), ZN => net136198);
   U9 : INV_X1 port map( A => b(2), ZN => net125371);
   U10 : NOR2_X1 port map( A1 => net153327, A2 => b(2), ZN => sel(0));
   U11 : AND3_X1 port map( A1 => b(2), A2 => n2, A3 => net136198, ZN => sel(2))
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BOOTHMUL is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL;

architecture SYN_MIXED of BOOTHMUL is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_DW01_sub_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   component MUX_5TO1_NBIT64_1
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_1
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_2
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_2
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_3
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_3
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_4
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_4
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_5
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_5
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_6
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_6
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_7
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_7
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_8
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_8
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_9
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_9
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_10
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_10
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_11
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_11
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_12
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_12
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_13
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_13
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_14
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_14
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_15
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component RCA_NBIT64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BE_BLOCK_15
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component MUX_5TO1_NBIT64_0
      port( A0, A1, A2, A3, A4 : in std_logic_vector (63 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto
            0));
   end component;
   
   component BE_BLOCK_0
      port( b : in std_logic_vector (2 downto 0);  sel : out std_logic_vector 
            (2 downto 0));
   end component;
   
   signal X_Logic0_port, selVector_15_2_port, selVector_15_1_port, 
      selVector_15_0_port, selVector_14_2_port, selVector_14_1_port, 
      selVector_14_0_port, selVector_13_2_port, selVector_13_1_port, 
      selVector_13_0_port, selVector_12_2_port, selVector_12_1_port, 
      selVector_12_0_port, selVector_11_2_port, selVector_11_1_port, 
      selVector_11_0_port, selVector_10_2_port, selVector_10_1_port, 
      selVector_10_0_port, selVector_9_2_port, selVector_9_1_port, 
      selVector_9_0_port, selVector_8_2_port, selVector_8_1_port, 
      selVector_8_0_port, selVector_7_2_port, selVector_7_1_port, 
      selVector_7_0_port, selVector_6_2_port, selVector_6_1_port, 
      selVector_6_0_port, selVector_5_2_port, selVector_5_1_port, 
      selVector_5_0_port, selVector_4_2_port, selVector_4_1_port, 
      selVector_4_0_port, selVector_3_2_port, selVector_3_1_port, 
      selVector_3_0_port, selVector_2_2_port, selVector_2_1_port, 
      selVector_2_0_port, selVector_1_2_port, selVector_1_1_port, 
      selVector_1_0_port, selVector_0_2_port, selVector_0_1_port, 
      selVector_0_0_port, muxOutVector_7_63_port, muxOutVector_7_62_port, 
      muxOutVector_7_61_port, muxOutVector_7_60_port, muxOutVector_7_59_port, 
      muxOutVector_7_58_port, muxOutVector_7_57_port, muxOutVector_7_56_port, 
      muxOutVector_7_55_port, muxOutVector_7_54_port, muxOutVector_7_53_port, 
      muxOutVector_7_52_port, muxOutVector_7_51_port, muxOutVector_7_50_port, 
      muxOutVector_7_49_port, muxOutVector_7_48_port, muxOutVector_7_47_port, 
      muxOutVector_7_46_port, muxOutVector_7_45_port, muxOutVector_7_44_port, 
      muxOutVector_7_43_port, muxOutVector_7_42_port, muxOutVector_7_41_port, 
      muxOutVector_7_40_port, muxOutVector_7_39_port, muxOutVector_7_38_port, 
      muxOutVector_7_37_port, muxOutVector_7_36_port, muxOutVector_7_35_port, 
      muxOutVector_7_34_port, muxOutVector_7_33_port, muxOutVector_7_32_port, 
      muxOutVector_7_31_port, muxOutVector_7_30_port, muxOutVector_7_29_port, 
      muxOutVector_7_28_port, muxOutVector_7_27_port, muxOutVector_7_26_port, 
      muxOutVector_7_25_port, muxOutVector_7_24_port, muxOutVector_7_23_port, 
      muxOutVector_7_22_port, muxOutVector_7_21_port, muxOutVector_7_20_port, 
      muxOutVector_7_19_port, muxOutVector_7_18_port, muxOutVector_7_17_port, 
      muxOutVector_7_16_port, muxOutVector_7_15_port, muxOutVector_7_14_port, 
      muxOutVector_7_13_port, muxOutVector_7_12_port, muxOutVector_7_11_port, 
      muxOutVector_7_10_port, muxOutVector_7_9_port, muxOutVector_7_8_port, 
      muxOutVector_7_7_port, muxOutVector_7_6_port, muxOutVector_7_5_port, 
      muxOutVector_7_4_port, muxOutVector_7_3_port, muxOutVector_7_2_port, 
      muxOutVector_7_1_port, muxOutVector_7_0_port, muxOutVector_6_63_port, 
      muxOutVector_6_62_port, muxOutVector_6_61_port, muxOutVector_6_60_port, 
      muxOutVector_6_59_port, muxOutVector_6_58_port, muxOutVector_6_57_port, 
      muxOutVector_6_56_port, muxOutVector_6_55_port, muxOutVector_6_54_port, 
      muxOutVector_6_53_port, muxOutVector_6_52_port, muxOutVector_6_51_port, 
      muxOutVector_6_50_port, muxOutVector_6_49_port, muxOutVector_6_48_port, 
      muxOutVector_6_47_port, muxOutVector_6_46_port, muxOutVector_6_45_port, 
      muxOutVector_6_44_port, muxOutVector_6_43_port, muxOutVector_6_42_port, 
      muxOutVector_6_41_port, muxOutVector_6_40_port, muxOutVector_6_39_port, 
      muxOutVector_6_38_port, muxOutVector_6_37_port, muxOutVector_6_36_port, 
      muxOutVector_6_35_port, muxOutVector_6_34_port, muxOutVector_6_33_port, 
      muxOutVector_6_32_port, muxOutVector_6_31_port, muxOutVector_6_30_port, 
      muxOutVector_6_29_port, muxOutVector_6_28_port, muxOutVector_6_27_port, 
      muxOutVector_6_26_port, muxOutVector_6_25_port, muxOutVector_6_24_port, 
      muxOutVector_6_23_port, muxOutVector_6_22_port, muxOutVector_6_21_port, 
      muxOutVector_6_20_port, muxOutVector_6_19_port, muxOutVector_6_18_port, 
      muxOutVector_6_17_port, muxOutVector_6_16_port, muxOutVector_6_15_port, 
      muxOutVector_6_14_port, muxOutVector_6_13_port, muxOutVector_6_12_port, 
      muxOutVector_6_11_port, muxOutVector_6_10_port, muxOutVector_6_9_port, 
      muxOutVector_6_8_port, muxOutVector_6_7_port, muxOutVector_6_6_port, 
      muxOutVector_6_5_port, muxOutVector_6_4_port, muxOutVector_6_3_port, 
      muxOutVector_6_2_port, muxOutVector_6_1_port, muxOutVector_6_0_port, 
      muxOutVector_5_63_port, muxOutVector_5_62_port, muxOutVector_5_61_port, 
      muxOutVector_5_60_port, muxOutVector_5_59_port, muxOutVector_5_58_port, 
      muxOutVector_5_57_port, muxOutVector_5_56_port, muxOutVector_5_55_port, 
      muxOutVector_5_54_port, muxOutVector_5_53_port, muxOutVector_5_52_port, 
      muxOutVector_5_51_port, muxOutVector_5_50_port, muxOutVector_5_49_port, 
      muxOutVector_5_48_port, muxOutVector_5_47_port, muxOutVector_5_46_port, 
      muxOutVector_5_45_port, muxOutVector_5_44_port, muxOutVector_5_43_port, 
      muxOutVector_5_42_port, muxOutVector_5_41_port, muxOutVector_5_40_port, 
      muxOutVector_5_39_port, muxOutVector_5_38_port, muxOutVector_5_37_port, 
      muxOutVector_5_36_port, muxOutVector_5_35_port, muxOutVector_5_34_port, 
      muxOutVector_5_33_port, muxOutVector_5_32_port, muxOutVector_5_31_port, 
      muxOutVector_5_30_port, muxOutVector_5_29_port, muxOutVector_5_28_port, 
      muxOutVector_5_27_port, muxOutVector_5_26_port, muxOutVector_5_25_port, 
      muxOutVector_5_24_port, muxOutVector_5_23_port, muxOutVector_5_22_port, 
      muxOutVector_5_21_port, muxOutVector_5_20_port, muxOutVector_5_19_port, 
      muxOutVector_5_18_port, muxOutVector_5_17_port, muxOutVector_5_16_port, 
      muxOutVector_5_15_port, muxOutVector_5_14_port, muxOutVector_5_13_port, 
      muxOutVector_5_12_port, muxOutVector_5_11_port, muxOutVector_5_10_port, 
      muxOutVector_5_9_port, muxOutVector_5_8_port, muxOutVector_5_7_port, 
      muxOutVector_5_6_port, muxOutVector_5_5_port, muxOutVector_5_4_port, 
      muxOutVector_5_3_port, muxOutVector_5_2_port, muxOutVector_5_1_port, 
      muxOutVector_5_0_port, muxOutVector_4_63_port, muxOutVector_4_62_port, 
      muxOutVector_4_61_port, muxOutVector_4_60_port, muxOutVector_4_59_port, 
      muxOutVector_4_58_port, muxOutVector_4_57_port, muxOutVector_4_56_port, 
      muxOutVector_4_55_port, muxOutVector_4_54_port, muxOutVector_4_53_port, 
      muxOutVector_4_52_port, muxOutVector_4_51_port, muxOutVector_4_50_port, 
      muxOutVector_4_49_port, muxOutVector_4_48_port, muxOutVector_4_47_port, 
      muxOutVector_4_46_port, muxOutVector_4_45_port, muxOutVector_4_44_port, 
      muxOutVector_4_43_port, muxOutVector_4_42_port, muxOutVector_4_41_port, 
      muxOutVector_4_40_port, muxOutVector_4_39_port, muxOutVector_4_38_port, 
      muxOutVector_4_37_port, muxOutVector_4_36_port, muxOutVector_4_35_port, 
      muxOutVector_4_34_port, muxOutVector_4_33_port, muxOutVector_4_32_port, 
      muxOutVector_4_31_port, muxOutVector_4_30_port, muxOutVector_4_29_port, 
      muxOutVector_4_28_port, muxOutVector_4_27_port, muxOutVector_4_26_port, 
      muxOutVector_4_25_port, muxOutVector_4_24_port, muxOutVector_4_23_port, 
      muxOutVector_4_22_port, muxOutVector_4_21_port, muxOutVector_4_20_port, 
      muxOutVector_4_19_port, muxOutVector_4_18_port, muxOutVector_4_17_port, 
      muxOutVector_4_16_port, muxOutVector_4_15_port, muxOutVector_4_14_port, 
      muxOutVector_4_13_port, muxOutVector_4_12_port, muxOutVector_4_11_port, 
      muxOutVector_4_10_port, muxOutVector_4_9_port, muxOutVector_4_8_port, 
      muxOutVector_4_7_port, muxOutVector_4_6_port, muxOutVector_4_5_port, 
      muxOutVector_4_4_port, muxOutVector_4_3_port, muxOutVector_4_2_port, 
      muxOutVector_4_1_port, muxOutVector_4_0_port, muxOutVector_3_63_port, 
      muxOutVector_3_62_port, muxOutVector_3_61_port, muxOutVector_3_60_port, 
      muxOutVector_3_59_port, muxOutVector_3_58_port, muxOutVector_3_57_port, 
      muxOutVector_3_56_port, muxOutVector_3_55_port, muxOutVector_3_54_port, 
      muxOutVector_3_53_port, muxOutVector_3_52_port, muxOutVector_3_51_port, 
      muxOutVector_3_50_port, muxOutVector_3_49_port, muxOutVector_3_48_port, 
      muxOutVector_3_47_port, muxOutVector_3_46_port, muxOutVector_3_45_port, 
      muxOutVector_3_44_port, muxOutVector_3_43_port, muxOutVector_3_42_port, 
      muxOutVector_3_41_port, muxOutVector_3_40_port, muxOutVector_3_39_port, 
      muxOutVector_3_38_port, muxOutVector_3_37_port, muxOutVector_3_36_port, 
      muxOutVector_3_35_port, muxOutVector_3_34_port, muxOutVector_3_33_port, 
      muxOutVector_3_32_port, muxOutVector_3_31_port, muxOutVector_3_30_port, 
      muxOutVector_3_29_port, muxOutVector_3_28_port, muxOutVector_3_27_port, 
      muxOutVector_3_26_port, muxOutVector_3_25_port, muxOutVector_3_24_port, 
      muxOutVector_3_23_port, muxOutVector_3_22_port, muxOutVector_3_21_port, 
      muxOutVector_3_20_port, muxOutVector_3_19_port, muxOutVector_3_18_port, 
      muxOutVector_3_17_port, muxOutVector_3_16_port, muxOutVector_3_15_port, 
      muxOutVector_3_14_port, muxOutVector_3_13_port, muxOutVector_3_12_port, 
      muxOutVector_3_11_port, muxOutVector_3_10_port, muxOutVector_3_9_port, 
      muxOutVector_3_8_port, muxOutVector_3_7_port, muxOutVector_3_6_port, 
      muxOutVector_3_5_port, muxOutVector_3_4_port, muxOutVector_3_3_port, 
      muxOutVector_3_2_port, muxOutVector_3_1_port, muxOutVector_3_0_port, 
      muxOutVector_2_63_port, muxOutVector_2_62_port, muxOutVector_2_61_port, 
      muxOutVector_2_60_port, muxOutVector_2_59_port, muxOutVector_2_58_port, 
      muxOutVector_2_57_port, muxOutVector_2_56_port, muxOutVector_2_55_port, 
      muxOutVector_2_54_port, muxOutVector_2_53_port, muxOutVector_2_52_port, 
      muxOutVector_2_51_port, muxOutVector_2_50_port, muxOutVector_2_49_port, 
      muxOutVector_2_48_port, muxOutVector_2_47_port, muxOutVector_2_46_port, 
      muxOutVector_2_45_port, muxOutVector_2_44_port, muxOutVector_2_43_port, 
      muxOutVector_2_42_port, muxOutVector_2_41_port, muxOutVector_2_40_port, 
      muxOutVector_2_39_port, muxOutVector_2_38_port, muxOutVector_2_37_port, 
      muxOutVector_2_36_port, muxOutVector_2_35_port, muxOutVector_2_34_port, 
      muxOutVector_2_33_port, muxOutVector_2_32_port, muxOutVector_2_31_port, 
      muxOutVector_2_30_port, muxOutVector_2_29_port, muxOutVector_2_28_port, 
      muxOutVector_2_27_port, muxOutVector_2_26_port, muxOutVector_2_25_port, 
      muxOutVector_2_24_port, muxOutVector_2_23_port, muxOutVector_2_22_port, 
      muxOutVector_2_21_port, muxOutVector_2_20_port, muxOutVector_2_19_port, 
      muxOutVector_2_18_port, muxOutVector_2_17_port, muxOutVector_2_16_port, 
      muxOutVector_2_15_port, muxOutVector_2_14_port, muxOutVector_2_13_port, 
      muxOutVector_2_12_port, muxOutVector_2_11_port, muxOutVector_2_10_port, 
      muxOutVector_2_9_port, muxOutVector_2_8_port, muxOutVector_2_7_port, 
      muxOutVector_2_6_port, muxOutVector_2_5_port, muxOutVector_2_4_port, 
      muxOutVector_2_3_port, muxOutVector_2_2_port, muxOutVector_2_1_port, 
      muxOutVector_2_0_port, muxOutVector_1_63_port, muxOutVector_1_62_port, 
      muxOutVector_1_61_port, muxOutVector_1_60_port, muxOutVector_1_59_port, 
      muxOutVector_1_58_port, muxOutVector_1_57_port, muxOutVector_1_56_port, 
      muxOutVector_1_55_port, muxOutVector_1_54_port, muxOutVector_1_53_port, 
      muxOutVector_1_52_port, muxOutVector_1_51_port, muxOutVector_1_50_port, 
      muxOutVector_1_49_port, muxOutVector_1_48_port, muxOutVector_1_47_port, 
      muxOutVector_1_46_port, muxOutVector_1_45_port, muxOutVector_1_44_port, 
      muxOutVector_1_43_port, muxOutVector_1_42_port, muxOutVector_1_41_port, 
      muxOutVector_1_40_port, muxOutVector_1_39_port, muxOutVector_1_38_port, 
      muxOutVector_1_37_port, muxOutVector_1_36_port, muxOutVector_1_35_port, 
      muxOutVector_1_34_port, muxOutVector_1_33_port, muxOutVector_1_32_port, 
      muxOutVector_1_31_port, muxOutVector_1_30_port, muxOutVector_1_29_port, 
      muxOutVector_1_28_port, muxOutVector_1_27_port, muxOutVector_1_26_port, 
      muxOutVector_1_25_port, muxOutVector_1_24_port, muxOutVector_1_23_port, 
      muxOutVector_1_22_port, muxOutVector_1_21_port, muxOutVector_1_20_port, 
      muxOutVector_1_19_port, muxOutVector_1_18_port, muxOutVector_1_17_port, 
      muxOutVector_1_16_port, muxOutVector_1_15_port, muxOutVector_1_14_port, 
      muxOutVector_1_13_port, muxOutVector_1_12_port, muxOutVector_1_11_port, 
      muxOutVector_1_10_port, muxOutVector_1_9_port, muxOutVector_1_8_port, 
      muxOutVector_1_7_port, muxOutVector_1_6_port, muxOutVector_1_5_port, 
      muxOutVector_1_4_port, muxOutVector_1_3_port, muxOutVector_1_2_port, 
      muxOutVector_1_1_port, muxOutVector_1_0_port, muxOutVector_0_63_port, 
      muxOutVector_0_62_port, muxOutVector_0_61_port, muxOutVector_0_60_port, 
      muxOutVector_0_59_port, muxOutVector_0_58_port, muxOutVector_0_57_port, 
      muxOutVector_0_56_port, muxOutVector_0_55_port, muxOutVector_0_54_port, 
      muxOutVector_0_53_port, muxOutVector_0_52_port, muxOutVector_0_51_port, 
      muxOutVector_0_50_port, muxOutVector_0_49_port, muxOutVector_0_48_port, 
      muxOutVector_0_47_port, muxOutVector_0_46_port, muxOutVector_0_45_port, 
      muxOutVector_0_44_port, muxOutVector_0_43_port, muxOutVector_0_42_port, 
      muxOutVector_0_41_port, muxOutVector_0_40_port, muxOutVector_0_39_port, 
      muxOutVector_0_38_port, muxOutVector_0_37_port, muxOutVector_0_36_port, 
      muxOutVector_0_35_port, muxOutVector_0_34_port, muxOutVector_0_33_port, 
      muxOutVector_0_32_port, muxOutVector_0_31_port, muxOutVector_0_30_port, 
      muxOutVector_0_29_port, muxOutVector_0_28_port, muxOutVector_0_27_port, 
      muxOutVector_0_26_port, muxOutVector_0_25_port, muxOutVector_0_24_port, 
      muxOutVector_0_23_port, muxOutVector_0_22_port, muxOutVector_0_21_port, 
      muxOutVector_0_20_port, muxOutVector_0_19_port, muxOutVector_0_18_port, 
      muxOutVector_0_17_port, muxOutVector_0_16_port, muxOutVector_0_15_port, 
      muxOutVector_0_14_port, muxOutVector_0_13_port, muxOutVector_0_12_port, 
      muxOutVector_0_11_port, muxOutVector_0_10_port, muxOutVector_0_9_port, 
      muxOutVector_0_8_port, muxOutVector_0_7_port, muxOutVector_0_6_port, 
      muxOutVector_0_5_port, muxOutVector_0_4_port, muxOutVector_0_3_port, 
      muxOutVector_0_2_port, muxOutVector_0_1_port, muxOutVector_0_0_port, 
      sumVector_14_63_port, sumVector_14_62_port, sumVector_14_61_port, 
      sumVector_14_60_port, sumVector_14_59_port, sumVector_14_58_port, 
      sumVector_14_57_port, sumVector_14_56_port, sumVector_14_55_port, 
      sumVector_14_54_port, sumVector_14_53_port, sumVector_14_52_port, 
      sumVector_14_51_port, sumVector_14_50_port, sumVector_14_49_port, 
      sumVector_14_48_port, sumVector_14_47_port, sumVector_14_46_port, 
      sumVector_14_45_port, sumVector_14_44_port, sumVector_14_43_port, 
      sumVector_14_42_port, sumVector_14_41_port, sumVector_14_40_port, 
      sumVector_14_39_port, sumVector_14_38_port, sumVector_14_37_port, 
      sumVector_14_36_port, sumVector_14_35_port, sumVector_14_34_port, 
      sumVector_14_33_port, sumVector_14_32_port, sumVector_14_31_port, 
      sumVector_14_30_port, sumVector_14_29_port, sumVector_14_28_port, 
      sumVector_14_27_port, sumVector_14_26_port, sumVector_14_25_port, 
      sumVector_14_24_port, sumVector_14_23_port, sumVector_14_22_port, 
      sumVector_14_21_port, sumVector_14_20_port, sumVector_14_19_port, 
      sumVector_14_18_port, sumVector_14_17_port, sumVector_14_16_port, 
      sumVector_14_15_port, sumVector_14_14_port, sumVector_14_13_port, 
      sumVector_14_12_port, sumVector_14_11_port, sumVector_14_10_port, 
      sumVector_14_9_port, sumVector_14_8_port, sumVector_14_7_port, 
      sumVector_14_6_port, sumVector_14_5_port, sumVector_14_4_port, 
      sumVector_14_3_port, sumVector_14_2_port, sumVector_14_1_port, 
      sumVector_14_0_port, sumVector_13_63_port, sumVector_13_62_port, 
      sumVector_13_61_port, sumVector_13_60_port, sumVector_13_59_port, 
      sumVector_13_58_port, sumVector_13_57_port, sumVector_13_56_port, 
      sumVector_13_55_port, sumVector_13_54_port, sumVector_13_53_port, 
      sumVector_13_52_port, sumVector_13_51_port, sumVector_13_50_port, 
      sumVector_13_49_port, sumVector_13_48_port, sumVector_13_47_port, 
      sumVector_13_46_port, sumVector_13_45_port, sumVector_13_44_port, 
      sumVector_13_43_port, sumVector_13_42_port, sumVector_13_41_port, 
      sumVector_13_40_port, sumVector_13_39_port, sumVector_13_38_port, 
      sumVector_13_37_port, sumVector_13_36_port, sumVector_13_35_port, 
      sumVector_13_34_port, sumVector_13_33_port, sumVector_13_32_port, 
      sumVector_13_31_port, sumVector_13_30_port, sumVector_13_29_port, 
      sumVector_13_28_port, sumVector_13_27_port, sumVector_13_26_port, 
      sumVector_13_25_port, sumVector_13_24_port, sumVector_13_23_port, 
      sumVector_13_22_port, sumVector_13_21_port, sumVector_13_20_port, 
      sumVector_13_19_port, sumVector_13_18_port, sumVector_13_17_port, 
      sumVector_13_16_port, sumVector_13_15_port, sumVector_13_14_port, 
      sumVector_13_13_port, sumVector_13_12_port, sumVector_13_11_port, 
      sumVector_13_10_port, sumVector_13_9_port, sumVector_13_8_port, 
      sumVector_13_7_port, sumVector_13_6_port, sumVector_13_5_port, 
      sumVector_13_4_port, sumVector_13_3_port, sumVector_13_2_port, 
      sumVector_13_1_port, sumVector_13_0_port, sumVector_12_63_port, 
      sumVector_12_62_port, sumVector_12_61_port, sumVector_12_60_port, 
      sumVector_12_59_port, sumVector_12_58_port, sumVector_12_57_port, 
      sumVector_12_56_port, sumVector_12_55_port, sumVector_12_54_port, 
      sumVector_12_53_port, sumVector_12_52_port, sumVector_12_51_port, 
      sumVector_12_50_port, sumVector_12_49_port, sumVector_12_48_port, 
      sumVector_12_47_port, sumVector_12_46_port, sumVector_12_45_port, 
      sumVector_12_44_port, sumVector_12_43_port, sumVector_12_42_port, 
      sumVector_12_41_port, sumVector_12_40_port, sumVector_12_39_port, 
      sumVector_12_38_port, sumVector_12_37_port, sumVector_12_36_port, 
      sumVector_12_35_port, sumVector_12_34_port, sumVector_12_33_port, 
      sumVector_12_32_port, sumVector_12_31_port, sumVector_12_30_port, 
      sumVector_12_29_port, sumVector_12_28_port, sumVector_12_27_port, 
      sumVector_12_26_port, sumVector_12_25_port, sumVector_12_24_port, 
      sumVector_12_23_port, sumVector_12_22_port, sumVector_12_21_port, 
      sumVector_12_20_port, sumVector_12_19_port, sumVector_12_18_port, 
      sumVector_12_17_port, sumVector_12_16_port, sumVector_12_15_port, 
      sumVector_12_14_port, sumVector_12_13_port, sumVector_12_12_port, 
      sumVector_12_11_port, sumVector_12_10_port, sumVector_12_9_port, 
      sumVector_12_8_port, sumVector_12_7_port, sumVector_12_6_port, 
      sumVector_12_5_port, sumVector_12_4_port, sumVector_12_3_port, 
      sumVector_12_2_port, sumVector_12_1_port, sumVector_12_0_port, 
      sumVector_11_63_port, sumVector_11_62_port, sumVector_11_61_port, 
      sumVector_11_60_port, sumVector_11_59_port, sumVector_11_58_port, 
      sumVector_11_57_port, sumVector_11_56_port, sumVector_11_55_port, 
      sumVector_11_54_port, sumVector_11_53_port, sumVector_11_52_port, 
      sumVector_11_51_port, sumVector_11_50_port, sumVector_11_49_port, 
      sumVector_11_48_port, sumVector_11_47_port, sumVector_11_46_port, 
      sumVector_11_45_port, sumVector_11_44_port, sumVector_11_43_port, 
      sumVector_11_42_port, sumVector_11_41_port, sumVector_11_40_port, 
      sumVector_11_39_port, sumVector_11_38_port, sumVector_11_37_port, 
      sumVector_11_36_port, sumVector_11_35_port, sumVector_11_34_port, 
      sumVector_11_33_port, sumVector_11_32_port, sumVector_11_31_port, 
      sumVector_11_30_port, sumVector_11_29_port, sumVector_11_28_port, 
      sumVector_11_27_port, sumVector_11_26_port, sumVector_11_25_port, 
      sumVector_11_24_port, sumVector_11_23_port, sumVector_11_22_port, 
      sumVector_11_21_port, sumVector_11_20_port, sumVector_11_19_port, 
      sumVector_11_18_port, sumVector_11_17_port, sumVector_11_16_port, 
      sumVector_11_15_port, sumVector_11_14_port, sumVector_11_13_port, 
      sumVector_11_12_port, sumVector_11_11_port, sumVector_11_10_port, 
      sumVector_11_9_port, sumVector_11_8_port, sumVector_11_7_port, 
      sumVector_11_6_port, sumVector_11_5_port, sumVector_11_4_port, 
      sumVector_11_3_port, sumVector_11_2_port, sumVector_11_1_port, 
      sumVector_11_0_port, sumVector_10_63_port, sumVector_10_62_port, 
      sumVector_10_61_port, sumVector_10_60_port, sumVector_10_59_port, 
      sumVector_10_58_port, sumVector_10_57_port, sumVector_10_56_port, 
      sumVector_10_55_port, sumVector_10_54_port, sumVector_10_53_port, 
      sumVector_10_52_port, sumVector_10_51_port, sumVector_10_50_port, 
      sumVector_10_49_port, sumVector_10_48_port, sumVector_10_47_port, 
      sumVector_10_46_port, sumVector_10_45_port, sumVector_10_44_port, 
      sumVector_10_43_port, sumVector_10_42_port, sumVector_10_41_port, 
      sumVector_10_40_port, sumVector_10_39_port, sumVector_10_38_port, 
      sumVector_10_37_port, sumVector_10_36_port, sumVector_10_35_port, 
      sumVector_10_34_port, sumVector_10_33_port, sumVector_10_32_port, 
      sumVector_10_31_port, sumVector_10_30_port, sumVector_10_29_port, 
      sumVector_10_28_port, sumVector_10_27_port, sumVector_10_26_port, 
      sumVector_10_25_port, sumVector_10_24_port, sumVector_10_23_port, 
      sumVector_10_22_port, sumVector_10_21_port, sumVector_10_20_port, 
      sumVector_10_19_port, sumVector_10_18_port, sumVector_10_17_port, 
      sumVector_10_16_port, sumVector_10_15_port, sumVector_10_14_port, 
      sumVector_10_13_port, sumVector_10_12_port, sumVector_10_11_port, 
      sumVector_10_10_port, sumVector_10_9_port, sumVector_10_8_port, 
      sumVector_10_7_port, sumVector_10_6_port, sumVector_10_5_port, 
      sumVector_10_4_port, sumVector_10_3_port, sumVector_10_2_port, 
      sumVector_10_1_port, sumVector_10_0_port, sumVector_9_63_port, 
      sumVector_9_62_port, sumVector_9_61_port, sumVector_9_60_port, 
      sumVector_9_59_port, sumVector_9_58_port, sumVector_9_57_port, 
      sumVector_9_56_port, sumVector_9_55_port, sumVector_9_54_port, 
      sumVector_9_53_port, sumVector_9_52_port, sumVector_9_51_port, 
      sumVector_9_50_port, sumVector_9_49_port, sumVector_9_48_port, 
      sumVector_9_47_port, sumVector_9_46_port, sumVector_9_45_port, 
      sumVector_9_44_port, sumVector_9_43_port, sumVector_9_42_port, 
      sumVector_9_41_port, sumVector_9_40_port, sumVector_9_39_port, 
      sumVector_9_38_port, sumVector_9_37_port, sumVector_9_36_port, 
      sumVector_9_35_port, sumVector_9_34_port, sumVector_9_33_port, 
      sumVector_9_32_port, sumVector_9_31_port, sumVector_9_30_port, 
      sumVector_9_29_port, sumVector_9_28_port, sumVector_9_27_port, 
      sumVector_9_26_port, sumVector_9_25_port, sumVector_9_24_port, 
      sumVector_9_23_port, sumVector_9_22_port, sumVector_9_21_port, 
      sumVector_9_20_port, sumVector_9_19_port, sumVector_9_18_port, 
      sumVector_9_17_port, sumVector_9_16_port, sumVector_9_15_port, 
      sumVector_9_14_port, sumVector_9_13_port, sumVector_9_12_port, 
      sumVector_9_11_port, sumVector_9_10_port, sumVector_9_9_port, 
      sumVector_9_8_port, sumVector_9_7_port, sumVector_9_6_port, 
      sumVector_9_5_port, sumVector_9_4_port, sumVector_9_3_port, 
      sumVector_9_2_port, sumVector_9_1_port, sumVector_9_0_port, 
      sumVector_8_63_port, sumVector_8_62_port, sumVector_8_61_port, 
      sumVector_8_60_port, sumVector_8_59_port, sumVector_8_58_port, 
      sumVector_8_57_port, sumVector_8_56_port, sumVector_8_55_port, 
      sumVector_8_54_port, sumVector_8_53_port, sumVector_8_52_port, 
      sumVector_8_51_port, sumVector_8_50_port, sumVector_8_49_port, 
      sumVector_8_48_port, sumVector_8_47_port, sumVector_8_46_port, 
      sumVector_8_45_port, sumVector_8_44_port, sumVector_8_43_port, 
      sumVector_8_42_port, sumVector_8_41_port, sumVector_8_40_port, 
      sumVector_8_39_port, sumVector_8_38_port, sumVector_8_37_port, 
      sumVector_8_36_port, sumVector_8_35_port, sumVector_8_34_port, 
      sumVector_8_33_port, sumVector_8_32_port, sumVector_8_31_port, 
      sumVector_8_30_port, sumVector_8_29_port, sumVector_8_28_port, 
      sumVector_8_27_port, sumVector_8_26_port, sumVector_8_25_port, 
      sumVector_8_24_port, sumVector_8_23_port, sumVector_8_22_port, 
      sumVector_8_21_port, sumVector_8_20_port, sumVector_8_19_port, 
      sumVector_8_18_port, sumVector_8_17_port, sumVector_8_16_port, 
      sumVector_8_15_port, sumVector_8_14_port, sumVector_8_13_port, 
      sumVector_8_12_port, sumVector_8_11_port, sumVector_8_10_port, 
      sumVector_8_9_port, sumVector_8_8_port, sumVector_8_7_port, 
      sumVector_8_6_port, sumVector_8_5_port, sumVector_8_4_port, 
      sumVector_8_3_port, sumVector_8_2_port, sumVector_8_1_port, 
      sumVector_8_0_port, sumVector_7_63_port, sumVector_7_62_port, 
      sumVector_7_61_port, sumVector_7_60_port, sumVector_7_59_port, 
      sumVector_7_58_port, sumVector_7_57_port, sumVector_7_56_port, 
      sumVector_7_55_port, sumVector_7_54_port, sumVector_7_53_port, 
      sumVector_7_52_port, sumVector_7_51_port, sumVector_7_50_port, 
      sumVector_7_49_port, sumVector_7_48_port, sumVector_7_47_port, 
      sumVector_7_46_port, sumVector_7_45_port, sumVector_7_44_port, 
      sumVector_7_43_port, sumVector_7_42_port, sumVector_7_41_port, 
      sumVector_7_40_port, sumVector_7_39_port, sumVector_7_38_port, 
      sumVector_7_37_port, sumVector_7_36_port, sumVector_7_35_port, 
      sumVector_7_34_port, sumVector_7_33_port, sumVector_7_32_port, 
      sumVector_7_31_port, sumVector_7_30_port, sumVector_7_29_port, 
      sumVector_7_28_port, sumVector_7_27_port, sumVector_7_26_port, 
      sumVector_7_25_port, sumVector_7_24_port, sumVector_7_23_port, 
      sumVector_7_22_port, sumVector_7_21_port, sumVector_7_20_port, 
      sumVector_7_19_port, sumVector_7_18_port, sumVector_7_17_port, 
      sumVector_7_16_port, sumVector_7_15_port, sumVector_7_14_port, 
      sumVector_7_13_port, sumVector_7_12_port, sumVector_7_11_port, 
      sumVector_7_10_port, sumVector_7_9_port, sumVector_7_8_port, 
      sumVector_7_7_port, sumVector_7_6_port, sumVector_7_5_port, 
      sumVector_7_4_port, sumVector_7_3_port, sumVector_7_2_port, 
      sumVector_7_1_port, sumVector_7_0_port, sumVector_6_63_port, 
      sumVector_6_62_port, sumVector_6_61_port, sumVector_6_60_port, 
      sumVector_6_59_port, sumVector_6_58_port, sumVector_6_57_port, 
      sumVector_6_56_port, sumVector_6_55_port, sumVector_6_54_port, 
      sumVector_6_53_port, sumVector_6_52_port, sumVector_6_51_port, 
      sumVector_6_50_port, sumVector_6_49_port, sumVector_6_48_port, 
      sumVector_6_47_port, sumVector_6_46_port, sumVector_6_45_port, 
      sumVector_6_44_port, sumVector_6_43_port, sumVector_6_42_port, 
      sumVector_6_41_port, sumVector_6_40_port, sumVector_6_39_port, 
      sumVector_6_38_port, sumVector_6_37_port, sumVector_6_36_port, 
      sumVector_6_35_port, sumVector_6_34_port, sumVector_6_33_port, 
      sumVector_6_32_port, sumVector_6_31_port, sumVector_6_30_port, 
      sumVector_6_29_port, sumVector_6_28_port, sumVector_6_27_port, 
      sumVector_6_26_port, sumVector_6_25_port, sumVector_6_24_port, 
      sumVector_6_23_port, sumVector_6_22_port, sumVector_6_21_port, 
      sumVector_6_20_port, sumVector_6_19_port, sumVector_6_18_port, 
      sumVector_6_17_port, sumVector_6_16_port, sumVector_6_15_port, 
      sumVector_6_14_port, sumVector_6_13_port, sumVector_6_12_port, 
      sumVector_6_11_port, sumVector_6_10_port, sumVector_6_9_port, 
      sumVector_6_8_port, sumVector_6_7_port, sumVector_6_6_port, 
      sumVector_6_5_port, sumVector_6_4_port, sumVector_6_3_port, 
      sumVector_6_2_port, sumVector_6_1_port, sumVector_6_0_port, 
      sumVector_5_63_port, sumVector_5_62_port, sumVector_5_61_port, 
      sumVector_5_60_port, sumVector_5_59_port, sumVector_5_58_port, 
      sumVector_5_57_port, sumVector_5_56_port, sumVector_5_55_port, 
      sumVector_5_54_port, sumVector_5_53_port, sumVector_5_52_port, 
      sumVector_5_51_port, sumVector_5_50_port, sumVector_5_49_port, 
      sumVector_5_48_port, sumVector_5_47_port, sumVector_5_46_port, 
      sumVector_5_45_port, sumVector_5_44_port, sumVector_5_43_port, 
      sumVector_5_42_port, sumVector_5_41_port, sumVector_5_40_port, 
      sumVector_5_39_port, sumVector_5_38_port, sumVector_5_37_port, 
      sumVector_5_36_port, sumVector_5_35_port, sumVector_5_34_port, 
      sumVector_5_33_port, sumVector_5_32_port, sumVector_5_31_port, 
      sumVector_5_30_port, sumVector_5_29_port, sumVector_5_28_port, 
      sumVector_5_27_port, sumVector_5_26_port, sumVector_5_25_port, 
      sumVector_5_24_port, sumVector_5_23_port, sumVector_5_22_port, 
      sumVector_5_21_port, sumVector_5_20_port, sumVector_5_19_port, 
      sumVector_5_18_port, sumVector_5_17_port, sumVector_5_16_port, 
      sumVector_5_15_port, sumVector_5_14_port, sumVector_5_13_port, 
      sumVector_5_12_port, sumVector_5_11_port, sumVector_5_10_port, 
      sumVector_5_9_port, sumVector_5_8_port, sumVector_5_7_port, 
      sumVector_5_6_port, sumVector_5_5_port, sumVector_5_4_port, 
      sumVector_5_3_port, sumVector_5_2_port, sumVector_5_1_port, 
      sumVector_5_0_port, sumVector_4_63_port, sumVector_4_62_port, 
      sumVector_4_61_port, sumVector_4_60_port, sumVector_4_59_port, 
      sumVector_4_58_port, sumVector_4_57_port, sumVector_4_56_port, 
      sumVector_4_55_port, sumVector_4_54_port, sumVector_4_53_port, 
      sumVector_4_52_port, sumVector_4_51_port, sumVector_4_50_port, 
      sumVector_4_49_port, sumVector_4_48_port, sumVector_4_47_port, 
      sumVector_4_46_port, sumVector_4_45_port, sumVector_4_44_port, 
      sumVector_4_43_port, sumVector_4_42_port, sumVector_4_41_port, 
      sumVector_4_40_port, sumVector_4_39_port, sumVector_4_38_port, 
      sumVector_4_37_port, sumVector_4_36_port, sumVector_4_35_port, 
      sumVector_4_34_port, sumVector_4_33_port, sumVector_4_32_port, 
      sumVector_4_31_port, sumVector_4_30_port, sumVector_4_29_port, 
      sumVector_4_28_port, sumVector_4_27_port, sumVector_4_26_port, 
      sumVector_4_25_port, sumVector_4_24_port, sumVector_4_23_port, 
      sumVector_4_22_port, sumVector_4_21_port, sumVector_4_20_port, 
      sumVector_4_19_port, sumVector_4_18_port, sumVector_4_17_port, 
      sumVector_4_16_port, sumVector_4_15_port, sumVector_4_14_port, 
      sumVector_4_13_port, sumVector_4_12_port, sumVector_4_11_port, 
      sumVector_4_10_port, sumVector_4_9_port, sumVector_4_8_port, 
      sumVector_4_7_port, sumVector_4_6_port, sumVector_4_5_port, 
      sumVector_4_4_port, sumVector_4_3_port, sumVector_4_2_port, 
      sumVector_4_1_port, sumVector_4_0_port, sumVector_3_63_port, 
      sumVector_3_62_port, sumVector_3_61_port, sumVector_3_60_port, 
      sumVector_3_59_port, sumVector_3_58_port, sumVector_3_57_port, 
      sumVector_3_56_port, sumVector_3_55_port, sumVector_3_54_port, 
      sumVector_3_53_port, sumVector_3_52_port, sumVector_3_51_port, 
      sumVector_3_50_port, sumVector_3_49_port, sumVector_3_48_port, 
      sumVector_3_47_port, sumVector_3_46_port, sumVector_3_45_port, 
      sumVector_3_44_port, sumVector_3_43_port, sumVector_3_42_port, 
      sumVector_3_41_port, sumVector_3_40_port, sumVector_3_39_port, 
      sumVector_3_38_port, sumVector_3_37_port, sumVector_3_36_port, 
      sumVector_3_35_port, sumVector_3_34_port, sumVector_3_33_port, 
      sumVector_3_32_port, sumVector_3_31_port, sumVector_3_30_port, 
      sumVector_3_29_port, sumVector_3_28_port, sumVector_3_27_port, 
      sumVector_3_26_port, sumVector_3_25_port, sumVector_3_24_port, 
      sumVector_3_23_port, sumVector_3_22_port, sumVector_3_21_port, 
      sumVector_3_20_port, sumVector_3_19_port, sumVector_3_18_port, 
      sumVector_3_17_port, sumVector_3_16_port, sumVector_3_15_port, 
      sumVector_3_14_port, sumVector_3_13_port, sumVector_3_12_port, 
      sumVector_3_11_port, sumVector_3_10_port, sumVector_3_9_port, 
      sumVector_3_8_port, sumVector_3_7_port, sumVector_3_6_port, 
      sumVector_3_5_port, sumVector_3_4_port, sumVector_3_3_port, 
      sumVector_3_2_port, sumVector_3_1_port, sumVector_3_0_port, 
      sumVector_2_63_port, sumVector_2_62_port, sumVector_2_61_port, 
      sumVector_2_60_port, sumVector_2_59_port, sumVector_2_58_port, 
      sumVector_2_57_port, sumVector_2_56_port, sumVector_2_55_port, 
      sumVector_2_54_port, sumVector_2_53_port, sumVector_2_52_port, 
      sumVector_2_51_port, sumVector_2_50_port, sumVector_2_49_port, 
      sumVector_2_48_port, sumVector_2_47_port, sumVector_2_46_port, 
      sumVector_2_45_port, sumVector_2_44_port, sumVector_2_43_port, 
      sumVector_2_42_port, sumVector_2_41_port, sumVector_2_40_port, 
      sumVector_2_39_port, sumVector_2_38_port, sumVector_2_37_port, 
      sumVector_2_36_port, sumVector_2_35_port, sumVector_2_34_port, 
      sumVector_2_33_port, sumVector_2_32_port, sumVector_2_31_port, 
      sumVector_2_30_port, sumVector_2_29_port, sumVector_2_28_port, 
      sumVector_2_27_port, sumVector_2_26_port, sumVector_2_25_port, 
      sumVector_2_24_port, sumVector_2_23_port, sumVector_2_22_port, 
      sumVector_2_21_port, sumVector_2_20_port, sumVector_2_19_port, 
      sumVector_2_18_port, sumVector_2_17_port, sumVector_2_16_port, 
      sumVector_2_15_port, sumVector_2_14_port, sumVector_2_13_port, 
      sumVector_2_12_port, sumVector_2_11_port, sumVector_2_10_port, 
      sumVector_2_9_port, sumVector_2_8_port, sumVector_2_7_port, 
      sumVector_2_6_port, sumVector_2_5_port, sumVector_2_4_port, 
      sumVector_2_3_port, sumVector_2_2_port, sumVector_2_1_port, 
      sumVector_2_0_port, sumVector_1_63_port, sumVector_1_62_port, 
      sumVector_1_61_port, sumVector_1_60_port, sumVector_1_59_port, 
      sumVector_1_58_port, sumVector_1_57_port, sumVector_1_56_port, 
      sumVector_1_55_port, sumVector_1_54_port, sumVector_1_53_port, 
      sumVector_1_52_port, sumVector_1_51_port, sumVector_1_50_port, 
      sumVector_1_49_port, sumVector_1_48_port, sumVector_1_47_port, 
      sumVector_1_46_port, sumVector_1_45_port, sumVector_1_44_port, 
      sumVector_1_43_port, sumVector_1_42_port, sumVector_1_41_port, 
      sumVector_1_40_port, sumVector_1_39_port, sumVector_1_38_port, 
      sumVector_1_37_port, sumVector_1_36_port, sumVector_1_35_port, 
      sumVector_1_34_port, sumVector_1_33_port, sumVector_1_32_port, 
      sumVector_1_31_port, sumVector_1_30_port, sumVector_1_29_port, 
      sumVector_1_28_port, sumVector_1_27_port, sumVector_1_26_port, 
      sumVector_1_25_port, sumVector_1_24_port, sumVector_1_23_port, 
      sumVector_1_22_port, sumVector_1_21_port, sumVector_1_20_port, 
      sumVector_1_19_port, sumVector_1_18_port, sumVector_1_17_port, 
      sumVector_1_16_port, sumVector_1_15_port, sumVector_1_14_port, 
      sumVector_1_13_port, sumVector_1_12_port, sumVector_1_11_port, 
      sumVector_1_10_port, sumVector_1_9_port, sumVector_1_8_port, 
      sumVector_1_7_port, sumVector_1_6_port, sumVector_1_5_port, 
      sumVector_1_4_port, sumVector_1_3_port, sumVector_1_2_port, 
      sumVector_1_1_port, sumVector_1_0_port, muxOutVector_15_63_port, 
      muxOutVector_15_62_port, muxOutVector_15_61_port, muxOutVector_15_60_port
      , muxOutVector_15_59_port, muxOutVector_15_58_port, 
      muxOutVector_15_57_port, muxOutVector_15_56_port, muxOutVector_15_55_port
      , muxOutVector_15_54_port, muxOutVector_15_53_port, 
      muxOutVector_15_52_port, muxOutVector_15_51_port, muxOutVector_15_50_port
      , muxOutVector_15_49_port, muxOutVector_15_48_port, 
      muxOutVector_15_47_port, muxOutVector_15_46_port, muxOutVector_15_45_port
      , muxOutVector_15_44_port, muxOutVector_15_43_port, 
      muxOutVector_15_42_port, muxOutVector_15_41_port, muxOutVector_15_40_port
      , muxOutVector_15_39_port, muxOutVector_15_38_port, 
      muxOutVector_15_37_port, muxOutVector_15_36_port, muxOutVector_15_35_port
      , muxOutVector_15_34_port, muxOutVector_15_33_port, 
      muxOutVector_15_32_port, muxOutVector_15_31_port, muxOutVector_15_30_port
      , muxOutVector_15_29_port, muxOutVector_15_28_port, 
      muxOutVector_15_27_port, muxOutVector_15_26_port, muxOutVector_15_25_port
      , muxOutVector_15_24_port, muxOutVector_15_23_port, 
      muxOutVector_15_22_port, muxOutVector_15_21_port, muxOutVector_15_20_port
      , muxOutVector_15_19_port, muxOutVector_15_18_port, 
      muxOutVector_15_17_port, muxOutVector_15_16_port, muxOutVector_15_15_port
      , muxOutVector_15_14_port, muxOutVector_15_13_port, 
      muxOutVector_15_12_port, muxOutVector_15_11_port, muxOutVector_15_10_port
      , muxOutVector_15_9_port, muxOutVector_15_8_port, muxOutVector_15_7_port,
      muxOutVector_15_6_port, muxOutVector_15_5_port, muxOutVector_15_4_port, 
      muxOutVector_15_3_port, muxOutVector_15_2_port, muxOutVector_15_1_port, 
      muxOutVector_15_0_port, muxOutVector_14_63_port, muxOutVector_14_62_port,
      muxOutVector_14_61_port, muxOutVector_14_60_port, muxOutVector_14_59_port
      , muxOutVector_14_58_port, muxOutVector_14_57_port, 
      muxOutVector_14_56_port, muxOutVector_14_55_port, muxOutVector_14_54_port
      , muxOutVector_14_53_port, muxOutVector_14_52_port, 
      muxOutVector_14_51_port, muxOutVector_14_50_port, muxOutVector_14_49_port
      , muxOutVector_14_48_port, muxOutVector_14_47_port, 
      muxOutVector_14_46_port, muxOutVector_14_45_port, muxOutVector_14_44_port
      , muxOutVector_14_43_port, muxOutVector_14_42_port, 
      muxOutVector_14_41_port, muxOutVector_14_40_port, muxOutVector_14_39_port
      , muxOutVector_14_38_port, muxOutVector_14_37_port, 
      muxOutVector_14_36_port, muxOutVector_14_35_port, muxOutVector_14_34_port
      , muxOutVector_14_33_port, muxOutVector_14_32_port, 
      muxOutVector_14_31_port, muxOutVector_14_30_port, muxOutVector_14_29_port
      , muxOutVector_14_28_port, muxOutVector_14_27_port, 
      muxOutVector_14_26_port, muxOutVector_14_25_port, muxOutVector_14_24_port
      , muxOutVector_14_23_port, muxOutVector_14_22_port, 
      muxOutVector_14_21_port, muxOutVector_14_20_port, muxOutVector_14_19_port
      , muxOutVector_14_18_port, muxOutVector_14_17_port, 
      muxOutVector_14_16_port, muxOutVector_14_15_port, muxOutVector_14_14_port
      , muxOutVector_14_13_port, muxOutVector_14_12_port, 
      muxOutVector_14_11_port, muxOutVector_14_10_port, muxOutVector_14_9_port,
      muxOutVector_14_8_port, muxOutVector_14_7_port, muxOutVector_14_6_port, 
      muxOutVector_14_5_port, muxOutVector_14_4_port, muxOutVector_14_3_port, 
      muxOutVector_14_2_port, muxOutVector_14_1_port, muxOutVector_14_0_port, 
      muxOutVector_13_63_port, muxOutVector_13_62_port, muxOutVector_13_61_port
      , muxOutVector_13_60_port, muxOutVector_13_59_port, 
      muxOutVector_13_58_port, muxOutVector_13_57_port, muxOutVector_13_56_port
      , muxOutVector_13_55_port, muxOutVector_13_54_port, 
      muxOutVector_13_53_port, muxOutVector_13_52_port, muxOutVector_13_51_port
      , muxOutVector_13_50_port, muxOutVector_13_49_port, 
      muxOutVector_13_48_port, muxOutVector_13_47_port, muxOutVector_13_46_port
      , muxOutVector_13_45_port, muxOutVector_13_44_port, 
      muxOutVector_13_43_port, muxOutVector_13_42_port, muxOutVector_13_41_port
      , muxOutVector_13_40_port, muxOutVector_13_39_port, 
      muxOutVector_13_38_port, muxOutVector_13_37_port, muxOutVector_13_36_port
      , muxOutVector_13_35_port, muxOutVector_13_34_port, 
      muxOutVector_13_33_port, muxOutVector_13_32_port, muxOutVector_13_31_port
      , muxOutVector_13_30_port, muxOutVector_13_29_port, 
      muxOutVector_13_28_port, muxOutVector_13_27_port, muxOutVector_13_26_port
      , muxOutVector_13_25_port, muxOutVector_13_24_port, 
      muxOutVector_13_23_port, muxOutVector_13_22_port, muxOutVector_13_21_port
      , muxOutVector_13_20_port, muxOutVector_13_19_port, 
      muxOutVector_13_18_port, muxOutVector_13_17_port, muxOutVector_13_16_port
      , muxOutVector_13_15_port, muxOutVector_13_14_port, 
      muxOutVector_13_13_port, muxOutVector_13_12_port, muxOutVector_13_11_port
      , muxOutVector_13_10_port, muxOutVector_13_9_port, muxOutVector_13_8_port
      , muxOutVector_13_7_port, muxOutVector_13_6_port, muxOutVector_13_5_port,
      muxOutVector_13_4_port, muxOutVector_13_3_port, muxOutVector_13_2_port, 
      muxOutVector_13_1_port, muxOutVector_13_0_port, muxOutVector_12_63_port, 
      muxOutVector_12_62_port, muxOutVector_12_61_port, muxOutVector_12_60_port
      , muxOutVector_12_59_port, muxOutVector_12_58_port, 
      muxOutVector_12_57_port, muxOutVector_12_56_port, muxOutVector_12_55_port
      , muxOutVector_12_54_port, muxOutVector_12_53_port, 
      muxOutVector_12_52_port, muxOutVector_12_51_port, muxOutVector_12_50_port
      , muxOutVector_12_49_port, muxOutVector_12_48_port, 
      muxOutVector_12_47_port, muxOutVector_12_46_port, muxOutVector_12_45_port
      , muxOutVector_12_44_port, muxOutVector_12_43_port, 
      muxOutVector_12_42_port, muxOutVector_12_41_port, muxOutVector_12_40_port
      , muxOutVector_12_39_port, muxOutVector_12_38_port, 
      muxOutVector_12_37_port, muxOutVector_12_36_port, muxOutVector_12_35_port
      , muxOutVector_12_34_port, muxOutVector_12_33_port, 
      muxOutVector_12_32_port, muxOutVector_12_31_port, muxOutVector_12_30_port
      , muxOutVector_12_29_port, muxOutVector_12_28_port, 
      muxOutVector_12_27_port, muxOutVector_12_26_port, muxOutVector_12_25_port
      , muxOutVector_12_24_port, muxOutVector_12_23_port, 
      muxOutVector_12_22_port, muxOutVector_12_21_port, muxOutVector_12_20_port
      , muxOutVector_12_19_port, muxOutVector_12_18_port, 
      muxOutVector_12_17_port, muxOutVector_12_16_port, muxOutVector_12_15_port
      , muxOutVector_12_14_port, muxOutVector_12_13_port, 
      muxOutVector_12_12_port, muxOutVector_12_11_port, muxOutVector_12_10_port
      , muxOutVector_12_9_port, muxOutVector_12_8_port, muxOutVector_12_7_port,
      muxOutVector_12_6_port, muxOutVector_12_5_port, muxOutVector_12_4_port, 
      muxOutVector_12_3_port, muxOutVector_12_2_port, muxOutVector_12_1_port, 
      muxOutVector_12_0_port, muxOutVector_11_63_port, muxOutVector_11_62_port,
      muxOutVector_11_61_port, muxOutVector_11_60_port, muxOutVector_11_59_port
      , muxOutVector_11_58_port, muxOutVector_11_57_port, 
      muxOutVector_11_56_port, muxOutVector_11_55_port, muxOutVector_11_54_port
      , muxOutVector_11_53_port, muxOutVector_11_52_port, 
      muxOutVector_11_51_port, muxOutVector_11_50_port, muxOutVector_11_49_port
      , muxOutVector_11_48_port, muxOutVector_11_47_port, 
      muxOutVector_11_46_port, muxOutVector_11_45_port, muxOutVector_11_44_port
      , muxOutVector_11_43_port, muxOutVector_11_42_port, 
      muxOutVector_11_41_port, muxOutVector_11_40_port, muxOutVector_11_39_port
      , muxOutVector_11_38_port, muxOutVector_11_37_port, 
      muxOutVector_11_36_port, muxOutVector_11_35_port, muxOutVector_11_34_port
      , muxOutVector_11_33_port, muxOutVector_11_32_port, 
      muxOutVector_11_31_port, muxOutVector_11_30_port, muxOutVector_11_29_port
      , muxOutVector_11_28_port, muxOutVector_11_27_port, 
      muxOutVector_11_26_port, muxOutVector_11_25_port, muxOutVector_11_24_port
      , muxOutVector_11_23_port, muxOutVector_11_22_port, 
      muxOutVector_11_21_port, muxOutVector_11_20_port, muxOutVector_11_19_port
      , muxOutVector_11_18_port, muxOutVector_11_17_port, 
      muxOutVector_11_16_port, muxOutVector_11_15_port, muxOutVector_11_14_port
      , muxOutVector_11_13_port, muxOutVector_11_12_port, 
      muxOutVector_11_11_port, muxOutVector_11_10_port, muxOutVector_11_9_port,
      muxOutVector_11_8_port, muxOutVector_11_7_port, muxOutVector_11_6_port, 
      muxOutVector_11_5_port, muxOutVector_11_4_port, muxOutVector_11_3_port, 
      muxOutVector_11_2_port, muxOutVector_11_1_port, muxOutVector_11_0_port, 
      muxOutVector_10_63_port, muxOutVector_10_62_port, muxOutVector_10_61_port
      , muxOutVector_10_60_port, muxOutVector_10_59_port, 
      muxOutVector_10_58_port, muxOutVector_10_57_port, muxOutVector_10_56_port
      , muxOutVector_10_55_port, muxOutVector_10_54_port, 
      muxOutVector_10_53_port, muxOutVector_10_52_port, muxOutVector_10_51_port
      , muxOutVector_10_50_port, muxOutVector_10_49_port, 
      muxOutVector_10_48_port, muxOutVector_10_47_port, muxOutVector_10_46_port
      , muxOutVector_10_45_port, muxOutVector_10_44_port, 
      muxOutVector_10_43_port, muxOutVector_10_42_port, muxOutVector_10_41_port
      , muxOutVector_10_40_port, muxOutVector_10_39_port, 
      muxOutVector_10_38_port, muxOutVector_10_37_port, muxOutVector_10_36_port
      , muxOutVector_10_35_port, muxOutVector_10_34_port, 
      muxOutVector_10_33_port, muxOutVector_10_32_port, muxOutVector_10_31_port
      , muxOutVector_10_30_port, muxOutVector_10_29_port, 
      muxOutVector_10_28_port, muxOutVector_10_27_port, muxOutVector_10_26_port
      , muxOutVector_10_25_port, muxOutVector_10_24_port, 
      muxOutVector_10_23_port, muxOutVector_10_22_port, muxOutVector_10_21_port
      , muxOutVector_10_20_port, muxOutVector_10_19_port, 
      muxOutVector_10_18_port, muxOutVector_10_17_port, muxOutVector_10_16_port
      , muxOutVector_10_15_port, muxOutVector_10_14_port, 
      muxOutVector_10_13_port, muxOutVector_10_12_port, muxOutVector_10_11_port
      , muxOutVector_10_10_port, muxOutVector_10_9_port, muxOutVector_10_8_port
      , muxOutVector_10_7_port, muxOutVector_10_6_port, muxOutVector_10_5_port,
      muxOutVector_10_4_port, muxOutVector_10_3_port, muxOutVector_10_2_port, 
      muxOutVector_10_1_port, muxOutVector_10_0_port, muxOutVector_9_63_port, 
      muxOutVector_9_62_port, muxOutVector_9_61_port, muxOutVector_9_60_port, 
      muxOutVector_9_59_port, muxOutVector_9_58_port, muxOutVector_9_57_port, 
      muxOutVector_9_56_port, muxOutVector_9_55_port, muxOutVector_9_54_port, 
      muxOutVector_9_53_port, muxOutVector_9_52_port, muxOutVector_9_51_port, 
      muxOutVector_9_50_port, muxOutVector_9_49_port, muxOutVector_9_48_port, 
      muxOutVector_9_47_port, muxOutVector_9_46_port, muxOutVector_9_45_port, 
      muxOutVector_9_44_port, muxOutVector_9_43_port, muxOutVector_9_42_port, 
      muxOutVector_9_41_port, muxOutVector_9_40_port, muxOutVector_9_39_port, 
      muxOutVector_9_38_port, muxOutVector_9_37_port, muxOutVector_9_36_port, 
      muxOutVector_9_35_port, muxOutVector_9_34_port, muxOutVector_9_33_port, 
      muxOutVector_9_32_port, muxOutVector_9_31_port, muxOutVector_9_30_port, 
      muxOutVector_9_29_port, muxOutVector_9_28_port, muxOutVector_9_27_port, 
      muxOutVector_9_26_port, muxOutVector_9_25_port, muxOutVector_9_24_port, 
      muxOutVector_9_23_port, muxOutVector_9_22_port, muxOutVector_9_21_port, 
      muxOutVector_9_20_port, muxOutVector_9_19_port, muxOutVector_9_18_port, 
      muxOutVector_9_17_port, muxOutVector_9_16_port, muxOutVector_9_15_port, 
      muxOutVector_9_14_port, muxOutVector_9_13_port, muxOutVector_9_12_port, 
      muxOutVector_9_11_port, muxOutVector_9_10_port, muxOutVector_9_9_port, 
      muxOutVector_9_8_port, muxOutVector_9_7_port, muxOutVector_9_6_port, 
      muxOutVector_9_5_port, muxOutVector_9_4_port, muxOutVector_9_3_port, 
      muxOutVector_9_2_port, muxOutVector_9_1_port, muxOutVector_9_0_port, 
      muxOutVector_8_63_port, muxOutVector_8_62_port, muxOutVector_8_61_port, 
      muxOutVector_8_60_port, muxOutVector_8_59_port, muxOutVector_8_58_port, 
      muxOutVector_8_57_port, muxOutVector_8_56_port, muxOutVector_8_55_port, 
      muxOutVector_8_54_port, muxOutVector_8_53_port, muxOutVector_8_52_port, 
      muxOutVector_8_51_port, muxOutVector_8_50_port, muxOutVector_8_49_port, 
      muxOutVector_8_48_port, muxOutVector_8_47_port, muxOutVector_8_46_port, 
      muxOutVector_8_45_port, muxOutVector_8_44_port, muxOutVector_8_43_port, 
      muxOutVector_8_42_port, muxOutVector_8_41_port, muxOutVector_8_40_port, 
      muxOutVector_8_39_port, muxOutVector_8_38_port, muxOutVector_8_37_port, 
      muxOutVector_8_36_port, muxOutVector_8_35_port, muxOutVector_8_34_port, 
      muxOutVector_8_33_port, muxOutVector_8_32_port, muxOutVector_8_31_port, 
      muxOutVector_8_30_port, muxOutVector_8_29_port, muxOutVector_8_28_port, 
      muxOutVector_8_27_port, muxOutVector_8_26_port, muxOutVector_8_25_port, 
      muxOutVector_8_24_port, muxOutVector_8_23_port, muxOutVector_8_22_port, 
      muxOutVector_8_21_port, muxOutVector_8_20_port, muxOutVector_8_19_port, 
      muxOutVector_8_18_port, muxOutVector_8_17_port, muxOutVector_8_16_port, 
      muxOutVector_8_15_port, muxOutVector_8_14_port, muxOutVector_8_13_port, 
      muxOutVector_8_12_port, muxOutVector_8_11_port, muxOutVector_8_10_port, 
      muxOutVector_8_9_port, muxOutVector_8_8_port, muxOutVector_8_7_port, 
      muxOutVector_8_6_port, muxOutVector_8_5_port, muxOutVector_8_4_port, 
      muxOutVector_8_3_port, muxOutVector_8_2_port, muxOutVector_8_1_port, 
      muxOutVector_8_0_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   n97 <= '0';
   n98 <= '0';
   eb_0 : BE_BLOCK_0 port map( b(2) => B(1), b(1) => B(0), b(0) => 
                           X_Logic0_port, sel(2) => selVector_0_2_port, sel(1) 
                           => selVector_0_1_port, sel(0) => selVector_0_0_port)
                           ;
   mux_0 : MUX_5TO1_NBIT64_0 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n122, A1(62) => n126, 
                           A1(61) => n126, A1(60) => n126, A1(59) => n126, 
                           A1(58) => n126, A1(57) => n126, A1(56) => n126, 
                           A1(55) => n126, A1(54) => n126, A1(53) => n126, 
                           A1(52) => n126, A1(51) => n125, A1(50) => n125, 
                           A1(49) => n125, A1(48) => n125, A1(47) => n125, 
                           A1(46) => n125, A1(45) => n125, A1(44) => n125, 
                           A1(43) => n125, A1(42) => n125, A1(41) => n125, 
                           A1(40) => n124, A1(39) => n124, A1(38) => n124, 
                           A1(37) => n124, A1(36) => n124, A1(35) => n124, 
                           A1(34) => n124, A1(33) => n124, A1(32) => n124, 
                           A1(31) => n124, A1(30) => n377, A1(29) => n370, 
                           A1(28) => n363, A1(27) => n356, A1(26) => n349, 
                           A1(25) => n342, A1(24) => n335, A1(23) => n328, 
                           A1(22) => n321, A1(21) => n314, A1(20) => n307, 
                           A1(19) => n300, A1(18) => n293, A1(17) => n286, 
                           A1(16) => n279, A1(15) => n272, A1(14) => n265, 
                           A1(13) => n258, A1(12) => n251, A1(11) => n244, 
                           A1(10) => n237, A1(9) => n230, A1(8) => n223, A1(7) 
                           => n216, A1(6) => n209, A1(5) => n202, A1(4) => n195
                           , A1(3) => n185, A1(2) => n178, A1(1) => n176, A1(0)
                           => A(0), A2(63) => n527, A2(62) => n527, A2(61) => 
                           n526, A2(60) => n526, A2(59) => n526, A2(58) => n526
                           , A2(57) => n526, A2(56) => n526, A2(55) => n526, 
                           A2(54) => n526, A2(53) => n526, A2(52) => n526, 
                           A2(51) => n526, A2(50) => n526, A2(49) => n525, 
                           A2(48) => n525, A2(47) => n525, A2(46) => n525, 
                           A2(45) => n525, A2(44) => n525, A2(43) => n525, 
                           A2(42) => n525, A2(41) => n525, A2(40) => n525, 
                           A2(39) => n525, A2(38) => n525, A2(37) => n524, 
                           A2(36) => n524, A2(35) => n524, A2(34) => n524, 
                           A2(33) => n524, A2(32) => n524, A2(31) => n493, 
                           A2(30) => n489, A2(29) => n485, A2(28) => n481, 
                           A2(27) => n477, A2(26) => n473, A2(25) => n469, 
                           A2(24) => n465, A2(23) => n461, A2(22) => n457, 
                           A2(21) => n453, A2(20) => n449, A2(19) => n445, 
                           A2(18) => n441, A2(17) => n437, A2(16) => n433, 
                           A2(15) => n430, A2(14) => n426, A2(13) => n423, 
                           A2(12) => n420, A2(11) => n416, A2(10) => n412, 
                           A2(9) => n409, A2(8) => n405, A2(7) => n401, A2(6) 
                           => n399, A2(5) => n395, A2(4) => n31, A2(3) => n32, 
                           A2(2) => n33, A2(1) => n383, A2(0) => n168, A3(63) 
                           => n144, A3(62) => n156, A3(61) => n139, A3(60) => 
                           n139, A3(59) => n139, A3(58) => n139, A3(57) => n139
                           , A3(56) => n139, A3(55) => n139, A3(54) => n139, 
                           A3(53) => n139, A3(52) => n139, A3(51) => n138, 
                           A3(50) => n138, A3(49) => n138, A3(48) => n138, 
                           A3(47) => n138, A3(46) => n138, A3(45) => n138, 
                           A3(44) => n138, A3(43) => n138, A3(42) => n138, 
                           A3(41) => n138, A3(40) => n138, A3(39) => n137, 
                           A3(38) => n137, A3(37) => n137, A3(36) => n142, 
                           A3(35) => n151, A3(34) => n151, A3(33) => n151, 
                           A3(32) => n151, A3(31) => n377, A3(30) => n370, 
                           A3(29) => n363, A3(28) => n356, A3(27) => n349, 
                           A3(26) => n342, A3(25) => n335, A3(24) => n328, 
                           A3(23) => n321, A3(22) => n314, A3(21) => n307, 
                           A3(20) => n300, A3(19) => n293, A3(18) => n286, 
                           A3(17) => n279, A3(16) => n272, A3(15) => n265, 
                           A3(14) => n258, A3(13) => n251, A3(12) => n244, 
                           A3(11) => n237, A3(10) => n230, A3(9) => n223, A3(8)
                           => n216, A3(7) => n209, A3(6) => n202, A3(5) => n195
                           , A3(4) => n185, A3(3) => n178, A3(2) => n175, A3(1)
                           => A(0), A3(0) => X_Logic0_port, A4(63) => n496, 
                           A4(62) => n510, A4(61) => n510, A4(60) => n509, 
                           A4(59) => n509, A4(58) => n509, A4(57) => n509, 
                           A4(56) => n509, A4(55) => n509, A4(54) => n509, 
                           A4(53) => n509, A4(52) => n509, A4(51) => n509, 
                           A4(50) => n509, A4(49) => n509, A4(48) => n508, 
                           A4(47) => n508, A4(46) => n508, A4(45) => n508, 
                           A4(44) => n508, A4(43) => n508, A4(42) => n508, 
                           A4(41) => n508, A4(40) => n508, A4(39) => n508, 
                           A4(38) => n508, A4(37) => n508, A4(36) => n507, 
                           A4(35) => n507, A4(34) => n507, A4(33) => n507, 
                           A4(32) => n492, A4(31) => n488, A4(30) => n484, 
                           A4(29) => n480, A4(28) => n476, A4(27) => n472, 
                           A4(26) => n468, A4(25) => n464, A4(24) => n460, 
                           A4(23) => n456, A4(22) => n452, A4(21) => n448, 
                           A4(20) => n444, A4(19) => n440, A4(18) => n436, 
                           A4(17) => n432, A4(16) => n429, A4(15) => n425, 
                           A4(14) => n422, A4(13) => n419, A4(12) => n415, 
                           A4(11) => n411, A4(10) => n408, A4(9) => n404, A4(8)
                           => n400, A4(7) => n105, A4(6) => n394, A4(5) => n391
                           , A4(4) => n388, A4(3) => n386, A4(2) => n384, A4(1)
                           => n167, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_0_2_port, sel(1) => selVector_0_1_port, 
                           sel(0) => selVector_0_0_port, O(63) => 
                           muxOutVector_0_63_port, O(62) => 
                           muxOutVector_0_62_port, O(61) => 
                           muxOutVector_0_61_port, O(60) => 
                           muxOutVector_0_60_port, O(59) => 
                           muxOutVector_0_59_port, O(58) => 
                           muxOutVector_0_58_port, O(57) => 
                           muxOutVector_0_57_port, O(56) => 
                           muxOutVector_0_56_port, O(55) => 
                           muxOutVector_0_55_port, O(54) => 
                           muxOutVector_0_54_port, O(53) => 
                           muxOutVector_0_53_port, O(52) => 
                           muxOutVector_0_52_port, O(51) => 
                           muxOutVector_0_51_port, O(50) => 
                           muxOutVector_0_50_port, O(49) => 
                           muxOutVector_0_49_port, O(48) => 
                           muxOutVector_0_48_port, O(47) => 
                           muxOutVector_0_47_port, O(46) => 
                           muxOutVector_0_46_port, O(45) => 
                           muxOutVector_0_45_port, O(44) => 
                           muxOutVector_0_44_port, O(43) => 
                           muxOutVector_0_43_port, O(42) => 
                           muxOutVector_0_42_port, O(41) => 
                           muxOutVector_0_41_port, O(40) => 
                           muxOutVector_0_40_port, O(39) => 
                           muxOutVector_0_39_port, O(38) => 
                           muxOutVector_0_38_port, O(37) => 
                           muxOutVector_0_37_port, O(36) => 
                           muxOutVector_0_36_port, O(35) => 
                           muxOutVector_0_35_port, O(34) => 
                           muxOutVector_0_34_port, O(33) => 
                           muxOutVector_0_33_port, O(32) => 
                           muxOutVector_0_32_port, O(31) => 
                           muxOutVector_0_31_port, O(30) => 
                           muxOutVector_0_30_port, O(29) => 
                           muxOutVector_0_29_port, O(28) => 
                           muxOutVector_0_28_port, O(27) => 
                           muxOutVector_0_27_port, O(26) => 
                           muxOutVector_0_26_port, O(25) => 
                           muxOutVector_0_25_port, O(24) => 
                           muxOutVector_0_24_port, O(23) => 
                           muxOutVector_0_23_port, O(22) => 
                           muxOutVector_0_22_port, O(21) => 
                           muxOutVector_0_21_port, O(20) => 
                           muxOutVector_0_20_port, O(19) => 
                           muxOutVector_0_19_port, O(18) => 
                           muxOutVector_0_18_port, O(17) => 
                           muxOutVector_0_17_port, O(16) => 
                           muxOutVector_0_16_port, O(15) => 
                           muxOutVector_0_15_port, O(14) => 
                           muxOutVector_0_14_port, O(13) => 
                           muxOutVector_0_13_port, O(12) => 
                           muxOutVector_0_12_port, O(11) => 
                           muxOutVector_0_11_port, O(10) => 
                           muxOutVector_0_10_port, O(9) => 
                           muxOutVector_0_9_port, O(8) => muxOutVector_0_8_port
                           , O(7) => muxOutVector_0_7_port, O(6) => 
                           muxOutVector_0_6_port, O(5) => muxOutVector_0_5_port
                           , O(4) => muxOutVector_0_4_port, O(3) => 
                           muxOutVector_0_3_port, O(2) => muxOutVector_0_2_port
                           , O(1) => muxOutVector_0_1_port, O(0) => 
                           muxOutVector_0_0_port);
   eb_1 : BE_BLOCK_15 port map( b(2) => B(3), b(1) => B(2), b(0) => B(1), 
                           sel(2) => selVector_1_2_port, sel(1) => 
                           selVector_1_1_port, sel(0) => selVector_1_0_port);
   sum_1 : RCA_NBIT64_0 port map( A(63) => muxOutVector_0_63_port, A(62) => 
                           muxOutVector_0_62_port, A(61) => 
                           muxOutVector_0_61_port, A(60) => 
                           muxOutVector_0_60_port, A(59) => 
                           muxOutVector_0_59_port, A(58) => 
                           muxOutVector_0_58_port, A(57) => 
                           muxOutVector_0_57_port, A(56) => 
                           muxOutVector_0_56_port, A(55) => 
                           muxOutVector_0_55_port, A(54) => 
                           muxOutVector_0_54_port, A(53) => 
                           muxOutVector_0_53_port, A(52) => 
                           muxOutVector_0_52_port, A(51) => 
                           muxOutVector_0_51_port, A(50) => 
                           muxOutVector_0_50_port, A(49) => 
                           muxOutVector_0_49_port, A(48) => 
                           muxOutVector_0_48_port, A(47) => 
                           muxOutVector_0_47_port, A(46) => 
                           muxOutVector_0_46_port, A(45) => 
                           muxOutVector_0_45_port, A(44) => 
                           muxOutVector_0_44_port, A(43) => 
                           muxOutVector_0_43_port, A(42) => 
                           muxOutVector_0_42_port, A(41) => 
                           muxOutVector_0_41_port, A(40) => 
                           muxOutVector_0_40_port, A(39) => 
                           muxOutVector_0_39_port, A(38) => 
                           muxOutVector_0_38_port, A(37) => 
                           muxOutVector_0_37_port, A(36) => 
                           muxOutVector_0_36_port, A(35) => 
                           muxOutVector_0_35_port, A(34) => 
                           muxOutVector_0_34_port, A(33) => 
                           muxOutVector_0_33_port, A(32) => 
                           muxOutVector_0_32_port, A(31) => 
                           muxOutVector_0_31_port, A(30) => 
                           muxOutVector_0_30_port, A(29) => 
                           muxOutVector_0_29_port, A(28) => 
                           muxOutVector_0_28_port, A(27) => 
                           muxOutVector_0_27_port, A(26) => 
                           muxOutVector_0_26_port, A(25) => 
                           muxOutVector_0_25_port, A(24) => 
                           muxOutVector_0_24_port, A(23) => 
                           muxOutVector_0_23_port, A(22) => 
                           muxOutVector_0_22_port, A(21) => 
                           muxOutVector_0_21_port, A(20) => 
                           muxOutVector_0_20_port, A(19) => 
                           muxOutVector_0_19_port, A(18) => 
                           muxOutVector_0_18_port, A(17) => 
                           muxOutVector_0_17_port, A(16) => 
                           muxOutVector_0_16_port, A(15) => 
                           muxOutVector_0_15_port, A(14) => 
                           muxOutVector_0_14_port, A(13) => 
                           muxOutVector_0_13_port, A(12) => 
                           muxOutVector_0_12_port, A(11) => 
                           muxOutVector_0_11_port, A(10) => 
                           muxOutVector_0_10_port, A(9) => 
                           muxOutVector_0_9_port, A(8) => muxOutVector_0_8_port
                           , A(7) => muxOutVector_0_7_port, A(6) => 
                           muxOutVector_0_6_port, A(5) => muxOutVector_0_5_port
                           , A(4) => muxOutVector_0_4_port, A(3) => 
                           muxOutVector_0_3_port, A(2) => muxOutVector_0_2_port
                           , A(1) => muxOutVector_0_1_port, A(0) => 
                           muxOutVector_0_0_port, B(63) => 
                           muxOutVector_1_63_port, B(62) => 
                           muxOutVector_1_62_port, B(61) => 
                           muxOutVector_1_61_port, B(60) => 
                           muxOutVector_1_60_port, B(59) => 
                           muxOutVector_1_59_port, B(58) => 
                           muxOutVector_1_58_port, B(57) => 
                           muxOutVector_1_57_port, B(56) => 
                           muxOutVector_1_56_port, B(55) => 
                           muxOutVector_1_55_port, B(54) => 
                           muxOutVector_1_54_port, B(53) => 
                           muxOutVector_1_53_port, B(52) => 
                           muxOutVector_1_52_port, B(51) => 
                           muxOutVector_1_51_port, B(50) => 
                           muxOutVector_1_50_port, B(49) => 
                           muxOutVector_1_49_port, B(48) => 
                           muxOutVector_1_48_port, B(47) => 
                           muxOutVector_1_47_port, B(46) => 
                           muxOutVector_1_46_port, B(45) => 
                           muxOutVector_1_45_port, B(44) => 
                           muxOutVector_1_44_port, B(43) => 
                           muxOutVector_1_43_port, B(42) => 
                           muxOutVector_1_42_port, B(41) => 
                           muxOutVector_1_41_port, B(40) => 
                           muxOutVector_1_40_port, B(39) => 
                           muxOutVector_1_39_port, B(38) => 
                           muxOutVector_1_38_port, B(37) => 
                           muxOutVector_1_37_port, B(36) => 
                           muxOutVector_1_36_port, B(35) => 
                           muxOutVector_1_35_port, B(34) => 
                           muxOutVector_1_34_port, B(33) => 
                           muxOutVector_1_33_port, B(32) => 
                           muxOutVector_1_32_port, B(31) => 
                           muxOutVector_1_31_port, B(30) => 
                           muxOutVector_1_30_port, B(29) => 
                           muxOutVector_1_29_port, B(28) => 
                           muxOutVector_1_28_port, B(27) => 
                           muxOutVector_1_27_port, B(26) => 
                           muxOutVector_1_26_port, B(25) => 
                           muxOutVector_1_25_port, B(24) => 
                           muxOutVector_1_24_port, B(23) => 
                           muxOutVector_1_23_port, B(22) => 
                           muxOutVector_1_22_port, B(21) => 
                           muxOutVector_1_21_port, B(20) => 
                           muxOutVector_1_20_port, B(19) => 
                           muxOutVector_1_19_port, B(18) => 
                           muxOutVector_1_18_port, B(17) => 
                           muxOutVector_1_17_port, B(16) => 
                           muxOutVector_1_16_port, B(15) => 
                           muxOutVector_1_15_port, B(14) => 
                           muxOutVector_1_14_port, B(13) => 
                           muxOutVector_1_13_port, B(12) => 
                           muxOutVector_1_12_port, B(11) => 
                           muxOutVector_1_11_port, B(10) => 
                           muxOutVector_1_10_port, B(9) => 
                           muxOutVector_1_9_port, B(8) => muxOutVector_1_8_port
                           , B(7) => muxOutVector_1_7_port, B(6) => 
                           muxOutVector_1_6_port, B(5) => muxOutVector_1_5_port
                           , B(4) => muxOutVector_1_4_port, B(3) => 
                           muxOutVector_1_3_port, B(2) => muxOutVector_1_2_port
                           , B(1) => muxOutVector_1_1_port, B(0) => 
                           muxOutVector_1_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_1_63_port, S(62) => sumVector_1_62_port, 
                           S(61) => sumVector_1_61_port, S(60) => 
                           sumVector_1_60_port, S(59) => sumVector_1_59_port, 
                           S(58) => sumVector_1_58_port, S(57) => 
                           sumVector_1_57_port, S(56) => sumVector_1_56_port, 
                           S(55) => sumVector_1_55_port, S(54) => 
                           sumVector_1_54_port, S(53) => sumVector_1_53_port, 
                           S(52) => sumVector_1_52_port, S(51) => 
                           sumVector_1_51_port, S(50) => sumVector_1_50_port, 
                           S(49) => sumVector_1_49_port, S(48) => 
                           sumVector_1_48_port, S(47) => sumVector_1_47_port, 
                           S(46) => sumVector_1_46_port, S(45) => 
                           sumVector_1_45_port, S(44) => sumVector_1_44_port, 
                           S(43) => sumVector_1_43_port, S(42) => 
                           sumVector_1_42_port, S(41) => sumVector_1_41_port, 
                           S(40) => sumVector_1_40_port, S(39) => 
                           sumVector_1_39_port, S(38) => sumVector_1_38_port, 
                           S(37) => sumVector_1_37_port, S(36) => 
                           sumVector_1_36_port, S(35) => sumVector_1_35_port, 
                           S(34) => sumVector_1_34_port, S(33) => 
                           sumVector_1_33_port, S(32) => sumVector_1_32_port, 
                           S(31) => sumVector_1_31_port, S(30) => 
                           sumVector_1_30_port, S(29) => sumVector_1_29_port, 
                           S(28) => sumVector_1_28_port, S(27) => 
                           sumVector_1_27_port, S(26) => sumVector_1_26_port, 
                           S(25) => sumVector_1_25_port, S(24) => 
                           sumVector_1_24_port, S(23) => sumVector_1_23_port, 
                           S(22) => sumVector_1_22_port, S(21) => 
                           sumVector_1_21_port, S(20) => sumVector_1_20_port, 
                           S(19) => sumVector_1_19_port, S(18) => 
                           sumVector_1_18_port, S(17) => sumVector_1_17_port, 
                           S(16) => sumVector_1_16_port, S(15) => 
                           sumVector_1_15_port, S(14) => sumVector_1_14_port, 
                           S(13) => sumVector_1_13_port, S(12) => 
                           sumVector_1_12_port, S(11) => sumVector_1_11_port, 
                           S(10) => sumVector_1_10_port, S(9) => 
                           sumVector_1_9_port, S(8) => sumVector_1_8_port, S(7)
                           => sumVector_1_7_port, S(6) => sumVector_1_6_port, 
                           S(5) => sumVector_1_5_port, S(4) => 
                           sumVector_1_4_port, S(3) => sumVector_1_3_port, S(2)
                           => sumVector_1_2_port, S(1) => sumVector_1_1_port, 
                           S(0) => sumVector_1_0_port, Co => n_1036);
   mux_1 : MUX_5TO1_NBIT64_15 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n145, A1(62) => n131, 
                           A1(61) => n131, A1(60) => n131, A1(59) => n131, 
                           A1(58) => n131, A1(57) => n131, A1(56) => n131, 
                           A1(55) => n130, A1(54) => n131, A1(53) => n130, 
                           A1(52) => n130, A1(51) => n130, A1(50) => n130, 
                           A1(49) => n131, A1(48) => n131, A1(47) => n131, 
                           A1(46) => n131, A1(45) => n130, A1(44) => n130, 
                           A1(43) => n131, A1(42) => n130, A1(41) => n130, 
                           A1(40) => n130, A1(39) => n130, A1(38) => n130, 
                           A1(37) => n130, A1(36) => n130, A1(35) => n130, 
                           A1(34) => n130, A1(33) => n130, A1(32) => n379, 
                           A1(31) => n372, A1(30) => n365, A1(29) => n358, 
                           A1(28) => n351, A1(27) => n344, A1(26) => n337, 
                           A1(25) => n330, A1(24) => n323, A1(23) => n316, 
                           A1(22) => n309, A1(21) => n302, A1(20) => n295, 
                           A1(19) => n288, A1(18) => n281, A1(17) => n274, 
                           A1(16) => n267, A1(15) => n260, A1(14) => n253, 
                           A1(13) => n246, A1(12) => n239, A1(11) => n232, 
                           A1(10) => n225, A1(9) => n218, A1(8) => n211, A1(7) 
                           => n204, A1(6) => n197, A1(5) => n185, A1(4) => n178
                           , A1(3) => n177, A1(2) => A(0), A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n519, A2(62) => n518, A2(61) => n519, A2(60) => n519
                           , A2(59) => n519, A2(58) => n519, A2(57) => n519, 
                           A2(56) => n520, A2(55) => n520, A2(54) => n520, 
                           A2(53) => n520, A2(52) => n521, A2(51) => n521, 
                           A2(50) => n521, A2(49) => n521, A2(48) => n521, 
                           A2(47) => n521, A2(46) => n521, A2(45) => n522, 
                           A2(44) => n522, A2(43) => n522, A2(42) => n522, 
                           A2(41) => n522, A2(40) => n523, A2(39) => n523, 
                           A2(38) => n523, A2(37) => n524, A2(36) => n524, 
                           A2(35) => n524, A2(34) => n524, A2(33) => n493, 
                           A2(32) => n489, A2(31) => n485, A2(30) => n481, 
                           A2(29) => n477, A2(28) => n473, A2(27) => n469, 
                           A2(26) => n465, A2(25) => n461, A2(24) => n457, 
                           A2(23) => n453, A2(22) => n449, A2(21) => n445, 
                           A2(20) => n441, A2(19) => n437, A2(18) => n433, 
                           A2(17) => n430, A2(16) => n426, A2(15) => n423, 
                           A2(14) => n420, A2(13) => n416, A2(12) => n412, 
                           A2(11) => n409, A2(10) => n405, A2(9) => n401, A2(8)
                           => n397, A2(7) => n396, A2(6) => n392, A2(5) => n389
                           , A2(4) => n387, A2(3) => n384, A2(2) => n35, A2(1) 
                           => X_Logic0_port, A2(0) => X_Logic0_port, A3(63) => 
                           n145, A3(62) => n146, A3(61) => n145, A3(60) => n146
                           , A3(59) => n145, A3(58) => n145, A3(57) => n145, 
                           A3(56) => n145, A3(55) => n146, A3(54) => n146, 
                           A3(53) => n145, A3(52) => n145, A3(51) => n145, 
                           A3(50) => n146, A3(49) => n145, A3(48) => n146, 
                           A3(47) => n145, A3(46) => n146, A3(45) => n146, 
                           A3(44) => n146, A3(43) => n146, A3(42) => n145, 
                           A3(41) => n146, A3(40) => n146, A3(39) => n146, 
                           A3(38) => n145, A3(37) => n146, A3(36) => n146, 
                           A3(35) => n146, A3(34) => n146, A3(33) => n379, 
                           A3(32) => n372, A3(31) => n365, A3(30) => n358, 
                           A3(29) => n351, A3(28) => n344, A3(27) => n337, 
                           A3(26) => n330, A3(25) => n323, A3(24) => n316, 
                           A3(23) => n309, A3(22) => n302, A3(21) => n295, 
                           A3(20) => n288, A3(19) => n281, A3(18) => n274, 
                           A3(17) => n267, A3(16) => n260, A3(15) => n253, 
                           A3(14) => n246, A3(13) => n239, A3(12) => n232, 
                           A3(11) => n225, A3(10) => n218, A3(9) => n211, A3(8)
                           => n204, A3(7) => n197, A3(6) => n170, A3(5) => n178
                           , A3(4) => n174, A3(3) => A(0), A3(2) => 
                           X_Logic0_port, A3(1) => X_Logic0_port, A3(0) => 
                           X_Logic0_port, A4(63) => n512, A4(62) => n512, 
                           A4(61) => n512, A4(60) => n512, A4(59) => n512, 
                           A4(58) => n512, A4(57) => n512, A4(56) => n513, 
                           A4(55) => n513, A4(54) => n513, A4(53) => n513, 
                           A4(52) => n513, A4(51) => n514, A4(50) => n514, 
                           A4(49) => n514, A4(48) => n514, A4(47) => n514, 
                           A4(46) => n514, A4(45) => n514, A4(44) => n514, 
                           A4(43) => n514, A4(42) => n514, A4(41) => n514, 
                           A4(40) => n515, A4(39) => n515, A4(38) => n515, 
                           A4(37) => n515, A4(36) => n515, A4(35) => n514, 
                           A4(34) => n492, A4(33) => n488, A4(32) => n484, 
                           A4(31) => n480, A4(30) => n476, A4(29) => n472, 
                           A4(28) => n468, A4(27) => n464, A4(26) => n460, 
                           A4(25) => n456, A4(24) => n452, A4(23) => n448, 
                           A4(22) => n444, A4(21) => n440, A4(20) => n436, 
                           A4(19) => n432, A4(18) => n429, A4(17) => n425, 
                           A4(16) => n422, A4(15) => n419, A4(14) => n415, 
                           A4(13) => n411, A4(12) => n408, A4(11) => n404, 
                           A4(10) => n400, A4(9) => n104, A4(8) => n394, A4(7) 
                           => n391, A4(6) => n100, A4(5) => n386, A4(4) => n383
                           , A4(3) => n35, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_1_2_port, sel(1) => selVector_1_1_port, 
                           sel(0) => selVector_1_0_port, O(63) => 
                           muxOutVector_1_63_port, O(62) => 
                           muxOutVector_1_62_port, O(61) => 
                           muxOutVector_1_61_port, O(60) => 
                           muxOutVector_1_60_port, O(59) => 
                           muxOutVector_1_59_port, O(58) => 
                           muxOutVector_1_58_port, O(57) => 
                           muxOutVector_1_57_port, O(56) => 
                           muxOutVector_1_56_port, O(55) => 
                           muxOutVector_1_55_port, O(54) => 
                           muxOutVector_1_54_port, O(53) => 
                           muxOutVector_1_53_port, O(52) => 
                           muxOutVector_1_52_port, O(51) => 
                           muxOutVector_1_51_port, O(50) => 
                           muxOutVector_1_50_port, O(49) => 
                           muxOutVector_1_49_port, O(48) => 
                           muxOutVector_1_48_port, O(47) => 
                           muxOutVector_1_47_port, O(46) => 
                           muxOutVector_1_46_port, O(45) => 
                           muxOutVector_1_45_port, O(44) => 
                           muxOutVector_1_44_port, O(43) => 
                           muxOutVector_1_43_port, O(42) => 
                           muxOutVector_1_42_port, O(41) => 
                           muxOutVector_1_41_port, O(40) => 
                           muxOutVector_1_40_port, O(39) => 
                           muxOutVector_1_39_port, O(38) => 
                           muxOutVector_1_38_port, O(37) => 
                           muxOutVector_1_37_port, O(36) => 
                           muxOutVector_1_36_port, O(35) => 
                           muxOutVector_1_35_port, O(34) => 
                           muxOutVector_1_34_port, O(33) => 
                           muxOutVector_1_33_port, O(32) => 
                           muxOutVector_1_32_port, O(31) => 
                           muxOutVector_1_31_port, O(30) => 
                           muxOutVector_1_30_port, O(29) => 
                           muxOutVector_1_29_port, O(28) => 
                           muxOutVector_1_28_port, O(27) => 
                           muxOutVector_1_27_port, O(26) => 
                           muxOutVector_1_26_port, O(25) => 
                           muxOutVector_1_25_port, O(24) => 
                           muxOutVector_1_24_port, O(23) => 
                           muxOutVector_1_23_port, O(22) => 
                           muxOutVector_1_22_port, O(21) => 
                           muxOutVector_1_21_port, O(20) => 
                           muxOutVector_1_20_port, O(19) => 
                           muxOutVector_1_19_port, O(18) => 
                           muxOutVector_1_18_port, O(17) => 
                           muxOutVector_1_17_port, O(16) => 
                           muxOutVector_1_16_port, O(15) => 
                           muxOutVector_1_15_port, O(14) => 
                           muxOutVector_1_14_port, O(13) => 
                           muxOutVector_1_13_port, O(12) => 
                           muxOutVector_1_12_port, O(11) => 
                           muxOutVector_1_11_port, O(10) => 
                           muxOutVector_1_10_port, O(9) => 
                           muxOutVector_1_9_port, O(8) => muxOutVector_1_8_port
                           , O(7) => muxOutVector_1_7_port, O(6) => 
                           muxOutVector_1_6_port, O(5) => muxOutVector_1_5_port
                           , O(4) => muxOutVector_1_4_port, O(3) => 
                           muxOutVector_1_3_port, O(2) => muxOutVector_1_2_port
                           , O(1) => muxOutVector_1_1_port, O(0) => 
                           muxOutVector_1_0_port);
   eb_2 : BE_BLOCK_14 port map( b(2) => B(5), b(1) => B(4), b(0) => B(3), 
                           sel(2) => selVector_2_2_port, sel(1) => 
                           selVector_2_1_port, sel(0) => selVector_2_0_port);
   sum_2 : RCA_NBIT64_14 port map( A(63) => muxOutVector_2_63_port, A(62) => 
                           muxOutVector_2_62_port, A(61) => 
                           muxOutVector_2_61_port, A(60) => 
                           muxOutVector_2_60_port, A(59) => 
                           muxOutVector_2_59_port, A(58) => 
                           muxOutVector_2_58_port, A(57) => 
                           muxOutVector_2_57_port, A(56) => 
                           muxOutVector_2_56_port, A(55) => 
                           muxOutVector_2_55_port, A(54) => 
                           muxOutVector_2_54_port, A(53) => 
                           muxOutVector_2_53_port, A(52) => 
                           muxOutVector_2_52_port, A(51) => 
                           muxOutVector_2_51_port, A(50) => 
                           muxOutVector_2_50_port, A(49) => 
                           muxOutVector_2_49_port, A(48) => 
                           muxOutVector_2_48_port, A(47) => 
                           muxOutVector_2_47_port, A(46) => 
                           muxOutVector_2_46_port, A(45) => 
                           muxOutVector_2_45_port, A(44) => 
                           muxOutVector_2_44_port, A(43) => 
                           muxOutVector_2_43_port, A(42) => 
                           muxOutVector_2_42_port, A(41) => 
                           muxOutVector_2_41_port, A(40) => 
                           muxOutVector_2_40_port, A(39) => 
                           muxOutVector_2_39_port, A(38) => 
                           muxOutVector_2_38_port, A(37) => 
                           muxOutVector_2_37_port, A(36) => 
                           muxOutVector_2_36_port, A(35) => 
                           muxOutVector_2_35_port, A(34) => 
                           muxOutVector_2_34_port, A(33) => 
                           muxOutVector_2_33_port, A(32) => 
                           muxOutVector_2_32_port, A(31) => 
                           muxOutVector_2_31_port, A(30) => 
                           muxOutVector_2_30_port, A(29) => 
                           muxOutVector_2_29_port, A(28) => 
                           muxOutVector_2_28_port, A(27) => 
                           muxOutVector_2_27_port, A(26) => 
                           muxOutVector_2_26_port, A(25) => 
                           muxOutVector_2_25_port, A(24) => 
                           muxOutVector_2_24_port, A(23) => 
                           muxOutVector_2_23_port, A(22) => 
                           muxOutVector_2_22_port, A(21) => 
                           muxOutVector_2_21_port, A(20) => 
                           muxOutVector_2_20_port, A(19) => 
                           muxOutVector_2_19_port, A(18) => 
                           muxOutVector_2_18_port, A(17) => 
                           muxOutVector_2_17_port, A(16) => 
                           muxOutVector_2_16_port, A(15) => 
                           muxOutVector_2_15_port, A(14) => 
                           muxOutVector_2_14_port, A(13) => 
                           muxOutVector_2_13_port, A(12) => 
                           muxOutVector_2_12_port, A(11) => 
                           muxOutVector_2_11_port, A(10) => 
                           muxOutVector_2_10_port, A(9) => 
                           muxOutVector_2_9_port, A(8) => muxOutVector_2_8_port
                           , A(7) => muxOutVector_2_7_port, A(6) => 
                           muxOutVector_2_6_port, A(5) => muxOutVector_2_5_port
                           , A(4) => muxOutVector_2_4_port, A(3) => 
                           muxOutVector_2_3_port, A(2) => muxOutVector_2_2_port
                           , A(1) => muxOutVector_2_1_port, A(0) => 
                           muxOutVector_2_0_port, B(63) => sumVector_1_63_port,
                           B(62) => sumVector_1_62_port, B(61) => 
                           sumVector_1_61_port, B(60) => sumVector_1_60_port, 
                           B(59) => sumVector_1_59_port, B(58) => 
                           sumVector_1_58_port, B(57) => sumVector_1_57_port, 
                           B(56) => sumVector_1_56_port, B(55) => 
                           sumVector_1_55_port, B(54) => sumVector_1_54_port, 
                           B(53) => sumVector_1_53_port, B(52) => 
                           sumVector_1_52_port, B(51) => sumVector_1_51_port, 
                           B(50) => sumVector_1_50_port, B(49) => 
                           sumVector_1_49_port, B(48) => sumVector_1_48_port, 
                           B(47) => sumVector_1_47_port, B(46) => 
                           sumVector_1_46_port, B(45) => sumVector_1_45_port, 
                           B(44) => sumVector_1_44_port, B(43) => 
                           sumVector_1_43_port, B(42) => sumVector_1_42_port, 
                           B(41) => sumVector_1_41_port, B(40) => 
                           sumVector_1_40_port, B(39) => sumVector_1_39_port, 
                           B(38) => sumVector_1_38_port, B(37) => 
                           sumVector_1_37_port, B(36) => sumVector_1_36_port, 
                           B(35) => sumVector_1_35_port, B(34) => 
                           sumVector_1_34_port, B(33) => sumVector_1_33_port, 
                           B(32) => sumVector_1_32_port, B(31) => 
                           sumVector_1_31_port, B(30) => sumVector_1_30_port, 
                           B(29) => sumVector_1_29_port, B(28) => 
                           sumVector_1_28_port, B(27) => sumVector_1_27_port, 
                           B(26) => sumVector_1_26_port, B(25) => 
                           sumVector_1_25_port, B(24) => sumVector_1_24_port, 
                           B(23) => sumVector_1_23_port, B(22) => 
                           sumVector_1_22_port, B(21) => sumVector_1_21_port, 
                           B(20) => sumVector_1_20_port, B(19) => 
                           sumVector_1_19_port, B(18) => sumVector_1_18_port, 
                           B(17) => sumVector_1_17_port, B(16) => 
                           sumVector_1_16_port, B(15) => sumVector_1_15_port, 
                           B(14) => sumVector_1_14_port, B(13) => 
                           sumVector_1_13_port, B(12) => sumVector_1_12_port, 
                           B(11) => sumVector_1_11_port, B(10) => 
                           sumVector_1_10_port, B(9) => sumVector_1_9_port, 
                           B(8) => sumVector_1_8_port, B(7) => 
                           sumVector_1_7_port, B(6) => sumVector_1_6_port, B(5)
                           => sumVector_1_5_port, B(4) => sumVector_1_4_port, 
                           B(3) => sumVector_1_3_port, B(2) => 
                           sumVector_1_2_port, B(1) => sumVector_1_1_port, B(0)
                           => sumVector_1_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_2_63_port, S(62) => sumVector_2_62_port, 
                           S(61) => sumVector_2_61_port, S(60) => 
                           sumVector_2_60_port, S(59) => sumVector_2_59_port, 
                           S(58) => sumVector_2_58_port, S(57) => 
                           sumVector_2_57_port, S(56) => sumVector_2_56_port, 
                           S(55) => sumVector_2_55_port, S(54) => 
                           sumVector_2_54_port, S(53) => sumVector_2_53_port, 
                           S(52) => sumVector_2_52_port, S(51) => 
                           sumVector_2_51_port, S(50) => sumVector_2_50_port, 
                           S(49) => sumVector_2_49_port, S(48) => 
                           sumVector_2_48_port, S(47) => sumVector_2_47_port, 
                           S(46) => sumVector_2_46_port, S(45) => 
                           sumVector_2_45_port, S(44) => sumVector_2_44_port, 
                           S(43) => sumVector_2_43_port, S(42) => 
                           sumVector_2_42_port, S(41) => sumVector_2_41_port, 
                           S(40) => sumVector_2_40_port, S(39) => 
                           sumVector_2_39_port, S(38) => sumVector_2_38_port, 
                           S(37) => sumVector_2_37_port, S(36) => 
                           sumVector_2_36_port, S(35) => sumVector_2_35_port, 
                           S(34) => sumVector_2_34_port, S(33) => 
                           sumVector_2_33_port, S(32) => sumVector_2_32_port, 
                           S(31) => sumVector_2_31_port, S(30) => 
                           sumVector_2_30_port, S(29) => sumVector_2_29_port, 
                           S(28) => sumVector_2_28_port, S(27) => 
                           sumVector_2_27_port, S(26) => sumVector_2_26_port, 
                           S(25) => sumVector_2_25_port, S(24) => 
                           sumVector_2_24_port, S(23) => sumVector_2_23_port, 
                           S(22) => sumVector_2_22_port, S(21) => 
                           sumVector_2_21_port, S(20) => sumVector_2_20_port, 
                           S(19) => sumVector_2_19_port, S(18) => 
                           sumVector_2_18_port, S(17) => sumVector_2_17_port, 
                           S(16) => sumVector_2_16_port, S(15) => 
                           sumVector_2_15_port, S(14) => sumVector_2_14_port, 
                           S(13) => sumVector_2_13_port, S(12) => 
                           sumVector_2_12_port, S(11) => sumVector_2_11_port, 
                           S(10) => sumVector_2_10_port, S(9) => 
                           sumVector_2_9_port, S(8) => sumVector_2_8_port, S(7)
                           => sumVector_2_7_port, S(6) => sumVector_2_6_port, 
                           S(5) => sumVector_2_5_port, S(4) => 
                           sumVector_2_4_port, S(3) => sumVector_2_3_port, S(2)
                           => sumVector_2_2_port, S(1) => sumVector_2_1_port, 
                           S(0) => sumVector_2_0_port, Co => n_1037);
   mux_2 : MUX_5TO1_NBIT64_14 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n110, A1(62) => n110, 
                           A1(61) => n110, A1(60) => n111, A1(59) => n111, 
                           A1(58) => n111, A1(57) => n111, A1(56) => n111, 
                           A1(55) => n111, A1(54) => n111, A1(53) => n111, 
                           A1(52) => n111, A1(51) => n111, A1(50) => n113, 
                           A1(49) => n113, A1(48) => n113, A1(47) => n113, 
                           A1(46) => n113, A1(45) => n113, A1(44) => n114, 
                           A1(43) => n114, A1(42) => n113, A1(41) => n114, 
                           A1(40) => n114, A1(39) => n114, A1(38) => n114, 
                           A1(37) => n114, A1(36) => n114, A1(35) => n114, 
                           A1(34) => n378, A1(33) => n371, A1(32) => n364, 
                           A1(31) => n357, A1(30) => n350, A1(29) => n343, 
                           A1(28) => n336, A1(27) => n329, A1(26) => n322, 
                           A1(25) => n315, A1(24) => n308, A1(23) => n301, 
                           A1(22) => n294, A1(21) => n287, A1(20) => n280, 
                           A1(19) => n273, A1(18) => n266, A1(17) => n259, 
                           A1(16) => n252, A1(15) => n245, A1(14) => n238, 
                           A1(13) => n231, A1(12) => n224, A1(11) => n217, 
                           A1(10) => n210, A1(9) => n203, A1(8) => n196, A1(7) 
                           => n171, A1(6) => n172, A1(5) => n176, A1(4) => A(0)
                           , A1(3) => X_Logic0_port, A1(2) => X_Logic0_port, 
                           A1(1) => X_Logic0_port, A1(0) => X_Logic0_port, 
                           A2(63) => n533, A2(62) => n534, A2(61) => n534, 
                           A2(60) => n535, A2(59) => n535, A2(58) => n535, 
                           A2(57) => n535, A2(56) => n535, A2(55) => n535, 
                           A2(54) => n535, A2(53) => n535, A2(52) => n535, 
                           A2(51) => n535, A2(50) => n535, A2(49) => n535, 
                           A2(48) => n536, A2(47) => n536, A2(46) => n536, 
                           A2(45) => n537, A2(44) => n537, A2(43) => n537, 
                           A2(42) => n538, A2(41) => n538, A2(40) => n538, 
                           A2(39) => n538, A2(38) => n538, A2(37) => n538, 
                           A2(36) => n538, A2(35) => n494, A2(34) => n490, 
                           A2(33) => n486, A2(32) => n482, A2(31) => n478, 
                           A2(30) => n474, A2(29) => n470, A2(28) => n466, 
                           A2(27) => n462, A2(26) => n458, A2(25) => n454, 
                           A2(24) => n450, A2(23) => n446, A2(22) => n442, 
                           A2(21) => n438, A2(20) => n434, A2(19) => n431, 
                           A2(18) => n427, A2(17) => n424, A2(16) => n421, 
                           A2(15) => n417, A2(14) => n413, A2(13) => n410, 
                           A2(12) => n406, A2(11) => n402, A2(10) => n397, 
                           A2(9) => n396, A2(8) => n392, A2(7) => n388, A2(6) 
                           => n387, A2(5) => n383, A2(4) => n35, A2(3) => 
                           X_Logic0_port, A2(2) => X_Logic0_port, A2(1) => 
                           X_Logic0_port, A2(0) => X_Logic0_port, A3(63) => 
                           n143, A3(62) => n143, A3(61) => n144, A3(60) => n144
                           , A3(59) => n142, A3(58) => n143, A3(57) => n142, 
                           A3(56) => n142, A3(55) => n144, A3(54) => n144, 
                           A3(53) => n145, A3(52) => n144, A3(51) => n143, 
                           A3(50) => n143, A3(49) => n143, A3(48) => n142, 
                           A3(47) => n144, A3(46) => n143, A3(45) => n142, 
                           A3(44) => n142, A3(43) => n144, A3(42) => n143, 
                           A3(41) => n142, A3(40) => n142, A3(39) => n142, 
                           A3(38) => n142, A3(37) => n140, A3(36) => n140, 
                           A3(35) => n377, A3(34) => n370, A3(33) => n363, 
                           A3(32) => n356, A3(31) => n349, A3(30) => n342, 
                           A3(29) => n335, A3(28) => n328, A3(27) => n321, 
                           A3(26) => n314, A3(25) => n307, A3(24) => n300, 
                           A3(23) => n293, A3(22) => n286, A3(21) => n279, 
                           A3(20) => n272, A3(19) => n265, A3(18) => n258, 
                           A3(17) => n251, A3(16) => n244, A3(15) => n237, 
                           A3(14) => n230, A3(13) => n223, A3(12) => n216, 
                           A3(11) => n209, A3(10) => n202, A3(9) => n195, A3(8)
                           => n190, A3(7) => n173, A3(6) => n176, A3(5) => A(0)
                           , A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n512, A4(62) => 
                           n512, A4(61) => n515, A4(60) => n515, A4(59) => n515
                           , A4(58) => n516, A4(57) => n516, A4(56) => n516, 
                           A4(55) => n516, A4(54) => n516, A4(53) => n516, 
                           A4(52) => n516, A4(51) => n516, A4(50) => n516, 
                           A4(49) => n516, A4(48) => n517, A4(47) => n516, 
                           A4(46) => n510, A4(45) => n515, A4(44) => n515, 
                           A4(43) => n515, A4(42) => n512, A4(41) => n512, 
                           A4(40) => n512, A4(39) => n511, A4(38) => n511, 
                           A4(37) => n511, A4(36) => n492, A4(35) => n488, 
                           A4(34) => n484, A4(33) => n480, A4(32) => n476, 
                           A4(31) => n472, A4(30) => n468, A4(29) => n464, 
                           A4(28) => n460, A4(27) => n456, A4(26) => n452, 
                           A4(25) => n448, A4(24) => n444, A4(23) => n440, 
                           A4(22) => n436, A4(21) => n432, A4(20) => n429, 
                           A4(19) => n425, A4(18) => n422, A4(17) => n419, 
                           A4(16) => n415, A4(15) => n411, A4(14) => n408, 
                           A4(13) => n404, A4(12) => n400, A4(11) => n398, 
                           A4(10) => n394, A4(9) => n391, A4(8) => n100, A4(7) 
                           => n386, A4(6) => n99, A4(5) => n35, A4(4) => 
                           X_Logic0_port, A4(3) => X_Logic0_port, A4(2) => 
                           X_Logic0_port, A4(1) => X_Logic0_port, A4(0) => 
                           X_Logic0_port, sel(2) => selVector_2_2_port, sel(1) 
                           => selVector_2_1_port, sel(0) => selVector_2_0_port,
                           O(63) => muxOutVector_2_63_port, O(62) => 
                           muxOutVector_2_62_port, O(61) => 
                           muxOutVector_2_61_port, O(60) => 
                           muxOutVector_2_60_port, O(59) => 
                           muxOutVector_2_59_port, O(58) => 
                           muxOutVector_2_58_port, O(57) => 
                           muxOutVector_2_57_port, O(56) => 
                           muxOutVector_2_56_port, O(55) => 
                           muxOutVector_2_55_port, O(54) => 
                           muxOutVector_2_54_port, O(53) => 
                           muxOutVector_2_53_port, O(52) => 
                           muxOutVector_2_52_port, O(51) => 
                           muxOutVector_2_51_port, O(50) => 
                           muxOutVector_2_50_port, O(49) => 
                           muxOutVector_2_49_port, O(48) => 
                           muxOutVector_2_48_port, O(47) => 
                           muxOutVector_2_47_port, O(46) => 
                           muxOutVector_2_46_port, O(45) => 
                           muxOutVector_2_45_port, O(44) => 
                           muxOutVector_2_44_port, O(43) => 
                           muxOutVector_2_43_port, O(42) => 
                           muxOutVector_2_42_port, O(41) => 
                           muxOutVector_2_41_port, O(40) => 
                           muxOutVector_2_40_port, O(39) => 
                           muxOutVector_2_39_port, O(38) => 
                           muxOutVector_2_38_port, O(37) => 
                           muxOutVector_2_37_port, O(36) => 
                           muxOutVector_2_36_port, O(35) => 
                           muxOutVector_2_35_port, O(34) => 
                           muxOutVector_2_34_port, O(33) => 
                           muxOutVector_2_33_port, O(32) => 
                           muxOutVector_2_32_port, O(31) => 
                           muxOutVector_2_31_port, O(30) => 
                           muxOutVector_2_30_port, O(29) => 
                           muxOutVector_2_29_port, O(28) => 
                           muxOutVector_2_28_port, O(27) => 
                           muxOutVector_2_27_port, O(26) => 
                           muxOutVector_2_26_port, O(25) => 
                           muxOutVector_2_25_port, O(24) => 
                           muxOutVector_2_24_port, O(23) => 
                           muxOutVector_2_23_port, O(22) => 
                           muxOutVector_2_22_port, O(21) => 
                           muxOutVector_2_21_port, O(20) => 
                           muxOutVector_2_20_port, O(19) => 
                           muxOutVector_2_19_port, O(18) => 
                           muxOutVector_2_18_port, O(17) => 
                           muxOutVector_2_17_port, O(16) => 
                           muxOutVector_2_16_port, O(15) => 
                           muxOutVector_2_15_port, O(14) => 
                           muxOutVector_2_14_port, O(13) => 
                           muxOutVector_2_13_port, O(12) => 
                           muxOutVector_2_12_port, O(11) => 
                           muxOutVector_2_11_port, O(10) => 
                           muxOutVector_2_10_port, O(9) => 
                           muxOutVector_2_9_port, O(8) => muxOutVector_2_8_port
                           , O(7) => muxOutVector_2_7_port, O(6) => 
                           muxOutVector_2_6_port, O(5) => muxOutVector_2_5_port
                           , O(4) => muxOutVector_2_4_port, O(3) => 
                           muxOutVector_2_3_port, O(2) => muxOutVector_2_2_port
                           , O(1) => muxOutVector_2_1_port, O(0) => 
                           muxOutVector_2_0_port);
   eb_3 : BE_BLOCK_13 port map( b(2) => B(7), b(1) => B(6), b(0) => B(5), 
                           sel(2) => selVector_3_2_port, sel(1) => 
                           selVector_3_1_port, sel(0) => selVector_3_0_port);
   sum_3 : RCA_NBIT64_13 port map( A(63) => muxOutVector_3_63_port, A(62) => 
                           muxOutVector_3_62_port, A(61) => 
                           muxOutVector_3_61_port, A(60) => 
                           muxOutVector_3_60_port, A(59) => 
                           muxOutVector_3_59_port, A(58) => 
                           muxOutVector_3_58_port, A(57) => 
                           muxOutVector_3_57_port, A(56) => 
                           muxOutVector_3_56_port, A(55) => 
                           muxOutVector_3_55_port, A(54) => 
                           muxOutVector_3_54_port, A(53) => 
                           muxOutVector_3_53_port, A(52) => 
                           muxOutVector_3_52_port, A(51) => 
                           muxOutVector_3_51_port, A(50) => 
                           muxOutVector_3_50_port, A(49) => 
                           muxOutVector_3_49_port, A(48) => 
                           muxOutVector_3_48_port, A(47) => 
                           muxOutVector_3_47_port, A(46) => 
                           muxOutVector_3_46_port, A(45) => 
                           muxOutVector_3_45_port, A(44) => 
                           muxOutVector_3_44_port, A(43) => 
                           muxOutVector_3_43_port, A(42) => 
                           muxOutVector_3_42_port, A(41) => 
                           muxOutVector_3_41_port, A(40) => 
                           muxOutVector_3_40_port, A(39) => 
                           muxOutVector_3_39_port, A(38) => 
                           muxOutVector_3_38_port, A(37) => 
                           muxOutVector_3_37_port, A(36) => 
                           muxOutVector_3_36_port, A(35) => 
                           muxOutVector_3_35_port, A(34) => 
                           muxOutVector_3_34_port, A(33) => 
                           muxOutVector_3_33_port, A(32) => 
                           muxOutVector_3_32_port, A(31) => 
                           muxOutVector_3_31_port, A(30) => 
                           muxOutVector_3_30_port, A(29) => 
                           muxOutVector_3_29_port, A(28) => 
                           muxOutVector_3_28_port, A(27) => 
                           muxOutVector_3_27_port, A(26) => 
                           muxOutVector_3_26_port, A(25) => 
                           muxOutVector_3_25_port, A(24) => 
                           muxOutVector_3_24_port, A(23) => 
                           muxOutVector_3_23_port, A(22) => 
                           muxOutVector_3_22_port, A(21) => 
                           muxOutVector_3_21_port, A(20) => 
                           muxOutVector_3_20_port, A(19) => 
                           muxOutVector_3_19_port, A(18) => 
                           muxOutVector_3_18_port, A(17) => 
                           muxOutVector_3_17_port, A(16) => 
                           muxOutVector_3_16_port, A(15) => 
                           muxOutVector_3_15_port, A(14) => 
                           muxOutVector_3_14_port, A(13) => 
                           muxOutVector_3_13_port, A(12) => 
                           muxOutVector_3_12_port, A(11) => 
                           muxOutVector_3_11_port, A(10) => 
                           muxOutVector_3_10_port, A(9) => 
                           muxOutVector_3_9_port, A(8) => muxOutVector_3_8_port
                           , A(7) => muxOutVector_3_7_port, A(6) => 
                           muxOutVector_3_6_port, A(5) => muxOutVector_3_5_port
                           , A(4) => muxOutVector_3_4_port, A(3) => 
                           muxOutVector_3_3_port, A(2) => muxOutVector_3_2_port
                           , A(1) => muxOutVector_3_1_port, A(0) => 
                           muxOutVector_3_0_port, B(63) => sumVector_2_63_port,
                           B(62) => sumVector_2_62_port, B(61) => 
                           sumVector_2_61_port, B(60) => sumVector_2_60_port, 
                           B(59) => sumVector_2_59_port, B(58) => 
                           sumVector_2_58_port, B(57) => sumVector_2_57_port, 
                           B(56) => sumVector_2_56_port, B(55) => 
                           sumVector_2_55_port, B(54) => sumVector_2_54_port, 
                           B(53) => sumVector_2_53_port, B(52) => 
                           sumVector_2_52_port, B(51) => sumVector_2_51_port, 
                           B(50) => sumVector_2_50_port, B(49) => 
                           sumVector_2_49_port, B(48) => sumVector_2_48_port, 
                           B(47) => sumVector_2_47_port, B(46) => 
                           sumVector_2_46_port, B(45) => sumVector_2_45_port, 
                           B(44) => sumVector_2_44_port, B(43) => 
                           sumVector_2_43_port, B(42) => sumVector_2_42_port, 
                           B(41) => sumVector_2_41_port, B(40) => 
                           sumVector_2_40_port, B(39) => sumVector_2_39_port, 
                           B(38) => sumVector_2_38_port, B(37) => 
                           sumVector_2_37_port, B(36) => sumVector_2_36_port, 
                           B(35) => sumVector_2_35_port, B(34) => 
                           sumVector_2_34_port, B(33) => sumVector_2_33_port, 
                           B(32) => sumVector_2_32_port, B(31) => 
                           sumVector_2_31_port, B(30) => sumVector_2_30_port, 
                           B(29) => sumVector_2_29_port, B(28) => 
                           sumVector_2_28_port, B(27) => sumVector_2_27_port, 
                           B(26) => sumVector_2_26_port, B(25) => 
                           sumVector_2_25_port, B(24) => sumVector_2_24_port, 
                           B(23) => sumVector_2_23_port, B(22) => 
                           sumVector_2_22_port, B(21) => sumVector_2_21_port, 
                           B(20) => sumVector_2_20_port, B(19) => 
                           sumVector_2_19_port, B(18) => sumVector_2_18_port, 
                           B(17) => sumVector_2_17_port, B(16) => 
                           sumVector_2_16_port, B(15) => sumVector_2_15_port, 
                           B(14) => sumVector_2_14_port, B(13) => 
                           sumVector_2_13_port, B(12) => sumVector_2_12_port, 
                           B(11) => sumVector_2_11_port, B(10) => 
                           sumVector_2_10_port, B(9) => sumVector_2_9_port, 
                           B(8) => sumVector_2_8_port, B(7) => 
                           sumVector_2_7_port, B(6) => sumVector_2_6_port, B(5)
                           => sumVector_2_5_port, B(4) => sumVector_2_4_port, 
                           B(3) => sumVector_2_3_port, B(2) => 
                           sumVector_2_2_port, B(1) => sumVector_2_1_port, B(0)
                           => sumVector_2_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_3_63_port, S(62) => sumVector_3_62_port, 
                           S(61) => sumVector_3_61_port, S(60) => 
                           sumVector_3_60_port, S(59) => sumVector_3_59_port, 
                           S(58) => sumVector_3_58_port, S(57) => 
                           sumVector_3_57_port, S(56) => sumVector_3_56_port, 
                           S(55) => sumVector_3_55_port, S(54) => 
                           sumVector_3_54_port, S(53) => sumVector_3_53_port, 
                           S(52) => sumVector_3_52_port, S(51) => 
                           sumVector_3_51_port, S(50) => sumVector_3_50_port, 
                           S(49) => sumVector_3_49_port, S(48) => 
                           sumVector_3_48_port, S(47) => sumVector_3_47_port, 
                           S(46) => sumVector_3_46_port, S(45) => 
                           sumVector_3_45_port, S(44) => sumVector_3_44_port, 
                           S(43) => sumVector_3_43_port, S(42) => 
                           sumVector_3_42_port, S(41) => sumVector_3_41_port, 
                           S(40) => sumVector_3_40_port, S(39) => 
                           sumVector_3_39_port, S(38) => sumVector_3_38_port, 
                           S(37) => sumVector_3_37_port, S(36) => 
                           sumVector_3_36_port, S(35) => sumVector_3_35_port, 
                           S(34) => sumVector_3_34_port, S(33) => 
                           sumVector_3_33_port, S(32) => sumVector_3_32_port, 
                           S(31) => sumVector_3_31_port, S(30) => 
                           sumVector_3_30_port, S(29) => sumVector_3_29_port, 
                           S(28) => sumVector_3_28_port, S(27) => 
                           sumVector_3_27_port, S(26) => sumVector_3_26_port, 
                           S(25) => sumVector_3_25_port, S(24) => 
                           sumVector_3_24_port, S(23) => sumVector_3_23_port, 
                           S(22) => sumVector_3_22_port, S(21) => 
                           sumVector_3_21_port, S(20) => sumVector_3_20_port, 
                           S(19) => sumVector_3_19_port, S(18) => 
                           sumVector_3_18_port, S(17) => sumVector_3_17_port, 
                           S(16) => sumVector_3_16_port, S(15) => 
                           sumVector_3_15_port, S(14) => sumVector_3_14_port, 
                           S(13) => sumVector_3_13_port, S(12) => 
                           sumVector_3_12_port, S(11) => sumVector_3_11_port, 
                           S(10) => sumVector_3_10_port, S(9) => 
                           sumVector_3_9_port, S(8) => sumVector_3_8_port, S(7)
                           => sumVector_3_7_port, S(6) => sumVector_3_6_port, 
                           S(5) => sumVector_3_5_port, S(4) => 
                           sumVector_3_4_port, S(3) => sumVector_3_3_port, S(2)
                           => sumVector_3_2_port, S(1) => sumVector_3_1_port, 
                           S(0) => sumVector_3_0_port, Co => n_1038);
   mux_3 : MUX_5TO1_NBIT64_13 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n116, A1(62) => n127, 
                           A1(61) => n126, A1(60) => n127, A1(59) => n127, 
                           A1(58) => n127, A1(57) => n129, A1(56) => n129, 
                           A1(55) => n129, A1(54) => n129, A1(53) => n129, 
                           A1(52) => n129, A1(51) => n130, A1(50) => n128, 
                           A1(49) => n121, A1(48) => n106, A1(47) => n106, 
                           A1(46) => n106, A1(45) => n106, A1(44) => n106, 
                           A1(43) => n106, A1(42) => n106, A1(41) => n106, 
                           A1(40) => n106, A1(39) => n106, A1(38) => n106, 
                           A1(37) => n106, A1(36) => n378, A1(35) => n371, 
                           A1(34) => n364, A1(33) => n357, A1(32) => n350, 
                           A1(31) => n343, A1(30) => n336, A1(29) => n329, 
                           A1(28) => n322, A1(27) => n315, A1(26) => n308, 
                           A1(25) => n301, A1(24) => n294, A1(23) => n287, 
                           A1(22) => n280, A1(21) => n273, A1(20) => n266, 
                           A1(19) => n259, A1(18) => n252, A1(17) => n245, 
                           A1(16) => n238, A1(15) => n231, A1(14) => n224, 
                           A1(13) => n217, A1(12) => n210, A1(11) => n203, 
                           A1(10) => n196, A1(9) => n188, A1(8) => n184, A1(7) 
                           => n102, A1(6) => A(0), A1(5) => X_Logic0_port, 
                           A1(4) => X_Logic0_port, A1(3) => X_Logic0_port, 
                           A1(2) => X_Logic0_port, A1(1) => X_Logic0_port, 
                           A1(0) => X_Logic0_port, A2(63) => n518, A2(62) => 
                           n533, A2(61) => n527, A2(60) => n527, A2(59) => n527
                           , A2(58) => n527, A2(57) => n527, A2(56) => n527, 
                           A2(55) => n527, A2(54) => n527, A2(53) => n527, 
                           A2(52) => n527, A2(51) => n530, A2(50) => n530, 
                           A2(49) => n530, A2(48) => n530, A2(47) => n530, 
                           A2(46) => n530, A2(45) => n530, A2(44) => n530, 
                           A2(43) => n530, A2(42) => n530, A2(41) => n530, 
                           A2(40) => n530, A2(39) => n531, A2(38) => n531, 
                           A2(37) => n494, A2(36) => n490, A2(35) => n486, 
                           A2(34) => n482, A2(33) => n478, A2(32) => n474, 
                           A2(31) => n470, A2(30) => n466, A2(29) => n462, 
                           A2(28) => n458, A2(27) => n454, A2(26) => n450, 
                           A2(25) => n446, A2(24) => n442, A2(23) => n438, 
                           A2(22) => n434, A2(21) => n431, A2(20) => n427, 
                           A2(19) => n424, A2(18) => n421, A2(17) => n417, 
                           A2(16) => n413, A2(15) => n410, A2(14) => n406, 
                           A2(13) => n402, A2(12) => n105, A2(11) => n396, 
                           A2(10) => n392, A2(9) => n101, A2(8) => n387, A2(7) 
                           => n383, A2(6) => n169, A2(5) => X_Logic0_port, 
                           A2(4) => X_Logic0_port, A2(3) => X_Logic0_port, 
                           A2(2) => X_Logic0_port, A2(1) => X_Logic0_port, 
                           A2(0) => X_Logic0_port, A3(63) => n142, A3(62) => 
                           n141, A3(61) => n141, A3(60) => n141, A3(59) => n141
                           , A3(58) => n141, A3(57) => n141, A3(56) => n141, 
                           A3(55) => n141, A3(54) => n141, A3(53) => n141, 
                           A3(52) => n141, A3(51) => n141, A3(50) => n140, 
                           A3(49) => n140, A3(48) => n140, A3(47) => n140, 
                           A3(46) => n140, A3(45) => n140, A3(44) => n140, 
                           A3(43) => n140, A3(42) => n140, A3(41) => n140, 
                           A3(40) => n139, A3(39) => n139, A3(38) => n143, 
                           A3(37) => n375, A3(36) => n368, A3(35) => n361, 
                           A3(34) => n354, A3(33) => n347, A3(32) => n340, 
                           A3(31) => n333, A3(30) => n326, A3(29) => n319, 
                           A3(28) => n312, A3(27) => n305, A3(26) => n298, 
                           A3(25) => n291, A3(24) => n284, A3(23) => n277, 
                           A3(22) => n270, A3(21) => n263, A3(20) => n256, 
                           A3(19) => n249, A3(18) => n242, A3(17) => n235, 
                           A3(16) => n228, A3(15) => n221, A3(14) => n214, 
                           A3(13) => n207, A3(12) => n200, A3(11) => n193, 
                           A3(10) => n191, A3(9) => n183, A3(8) => n103, A3(7) 
                           => A(0), A3(6) => X_Logic0_port, A3(5) => 
                           X_Logic0_port, A3(4) => X_Logic0_port, A3(3) => 
                           X_Logic0_port, A3(2) => X_Logic0_port, A3(1) => 
                           X_Logic0_port, A3(0) => X_Logic0_port, A4(63) => 
                           n513, A4(62) => n513, A4(61) => n513, A4(60) => n513
                           , A4(59) => n513, A4(58) => n513, A4(57) => n513, 
                           A4(56) => n511, A4(55) => n511, A4(54) => n511, 
                           A4(53) => n511, A4(52) => n511, A4(51) => n511, 
                           A4(50) => n511, A4(49) => n511, A4(48) => n511, 
                           A4(47) => n510, A4(46) => n510, A4(45) => n510, 
                           A4(44) => n510, A4(43) => n510, A4(42) => n510, 
                           A4(41) => n510, A4(40) => n510, A4(39) => n510, 
                           A4(38) => n492, A4(37) => n488, A4(36) => n484, 
                           A4(35) => n480, A4(34) => n476, A4(33) => n472, 
                           A4(32) => n468, A4(31) => n464, A4(30) => n460, 
                           A4(29) => n456, A4(28) => n452, A4(27) => n448, 
                           A4(26) => n444, A4(25) => n440, A4(24) => n436, 
                           A4(23) => n432, A4(22) => n429, A4(21) => n425, 
                           A4(20) => n422, A4(19) => n419, A4(18) => n415, 
                           A4(17) => n411, A4(16) => n408, A4(15) => n404, 
                           A4(14) => n400, A4(13) => n104, A4(12) => n394, 
                           A4(11) => n391, A4(10) => n389, A4(9) => n386, A4(8)
                           => n99, A4(7) => n167, A4(6) => X_Logic0_port, A4(5)
                           => X_Logic0_port, A4(4) => X_Logic0_port, A4(3) => 
                           X_Logic0_port, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_3_2_port, sel(1) => selVector_3_1_port, 
                           sel(0) => selVector_3_0_port, O(63) => 
                           muxOutVector_3_63_port, O(62) => 
                           muxOutVector_3_62_port, O(61) => 
                           muxOutVector_3_61_port, O(60) => 
                           muxOutVector_3_60_port, O(59) => 
                           muxOutVector_3_59_port, O(58) => 
                           muxOutVector_3_58_port, O(57) => 
                           muxOutVector_3_57_port, O(56) => 
                           muxOutVector_3_56_port, O(55) => 
                           muxOutVector_3_55_port, O(54) => 
                           muxOutVector_3_54_port, O(53) => 
                           muxOutVector_3_53_port, O(52) => 
                           muxOutVector_3_52_port, O(51) => 
                           muxOutVector_3_51_port, O(50) => 
                           muxOutVector_3_50_port, O(49) => 
                           muxOutVector_3_49_port, O(48) => 
                           muxOutVector_3_48_port, O(47) => 
                           muxOutVector_3_47_port, O(46) => 
                           muxOutVector_3_46_port, O(45) => 
                           muxOutVector_3_45_port, O(44) => 
                           muxOutVector_3_44_port, O(43) => 
                           muxOutVector_3_43_port, O(42) => 
                           muxOutVector_3_42_port, O(41) => 
                           muxOutVector_3_41_port, O(40) => 
                           muxOutVector_3_40_port, O(39) => 
                           muxOutVector_3_39_port, O(38) => 
                           muxOutVector_3_38_port, O(37) => 
                           muxOutVector_3_37_port, O(36) => 
                           muxOutVector_3_36_port, O(35) => 
                           muxOutVector_3_35_port, O(34) => 
                           muxOutVector_3_34_port, O(33) => 
                           muxOutVector_3_33_port, O(32) => 
                           muxOutVector_3_32_port, O(31) => 
                           muxOutVector_3_31_port, O(30) => 
                           muxOutVector_3_30_port, O(29) => 
                           muxOutVector_3_29_port, O(28) => 
                           muxOutVector_3_28_port, O(27) => 
                           muxOutVector_3_27_port, O(26) => 
                           muxOutVector_3_26_port, O(25) => 
                           muxOutVector_3_25_port, O(24) => 
                           muxOutVector_3_24_port, O(23) => 
                           muxOutVector_3_23_port, O(22) => 
                           muxOutVector_3_22_port, O(21) => 
                           muxOutVector_3_21_port, O(20) => 
                           muxOutVector_3_20_port, O(19) => 
                           muxOutVector_3_19_port, O(18) => 
                           muxOutVector_3_18_port, O(17) => 
                           muxOutVector_3_17_port, O(16) => 
                           muxOutVector_3_16_port, O(15) => 
                           muxOutVector_3_15_port, O(14) => 
                           muxOutVector_3_14_port, O(13) => 
                           muxOutVector_3_13_port, O(12) => 
                           muxOutVector_3_12_port, O(11) => 
                           muxOutVector_3_11_port, O(10) => 
                           muxOutVector_3_10_port, O(9) => 
                           muxOutVector_3_9_port, O(8) => muxOutVector_3_8_port
                           , O(7) => muxOutVector_3_7_port, O(6) => 
                           muxOutVector_3_6_port, O(5) => muxOutVector_3_5_port
                           , O(4) => muxOutVector_3_4_port, O(3) => 
                           muxOutVector_3_3_port, O(2) => muxOutVector_3_2_port
                           , O(1) => muxOutVector_3_1_port, O(0) => 
                           muxOutVector_3_0_port);
   eb_4 : BE_BLOCK_12 port map( b(2) => B(9), b(1) => B(8), b(0) => B(7), 
                           sel(2) => selVector_4_2_port, sel(1) => 
                           selVector_4_1_port, sel(0) => selVector_4_0_port);
   sum_4 : RCA_NBIT64_12 port map( A(63) => muxOutVector_4_63_port, A(62) => 
                           muxOutVector_4_62_port, A(61) => 
                           muxOutVector_4_61_port, A(60) => 
                           muxOutVector_4_60_port, A(59) => 
                           muxOutVector_4_59_port, A(58) => 
                           muxOutVector_4_58_port, A(57) => 
                           muxOutVector_4_57_port, A(56) => 
                           muxOutVector_4_56_port, A(55) => 
                           muxOutVector_4_55_port, A(54) => 
                           muxOutVector_4_54_port, A(53) => 
                           muxOutVector_4_53_port, A(52) => 
                           muxOutVector_4_52_port, A(51) => 
                           muxOutVector_4_51_port, A(50) => 
                           muxOutVector_4_50_port, A(49) => 
                           muxOutVector_4_49_port, A(48) => 
                           muxOutVector_4_48_port, A(47) => 
                           muxOutVector_4_47_port, A(46) => 
                           muxOutVector_4_46_port, A(45) => 
                           muxOutVector_4_45_port, A(44) => 
                           muxOutVector_4_44_port, A(43) => 
                           muxOutVector_4_43_port, A(42) => 
                           muxOutVector_4_42_port, A(41) => 
                           muxOutVector_4_41_port, A(40) => 
                           muxOutVector_4_40_port, A(39) => 
                           muxOutVector_4_39_port, A(38) => 
                           muxOutVector_4_38_port, A(37) => 
                           muxOutVector_4_37_port, A(36) => 
                           muxOutVector_4_36_port, A(35) => 
                           muxOutVector_4_35_port, A(34) => 
                           muxOutVector_4_34_port, A(33) => 
                           muxOutVector_4_33_port, A(32) => 
                           muxOutVector_4_32_port, A(31) => 
                           muxOutVector_4_31_port, A(30) => 
                           muxOutVector_4_30_port, A(29) => 
                           muxOutVector_4_29_port, A(28) => 
                           muxOutVector_4_28_port, A(27) => 
                           muxOutVector_4_27_port, A(26) => 
                           muxOutVector_4_26_port, A(25) => 
                           muxOutVector_4_25_port, A(24) => 
                           muxOutVector_4_24_port, A(23) => 
                           muxOutVector_4_23_port, A(22) => 
                           muxOutVector_4_22_port, A(21) => 
                           muxOutVector_4_21_port, A(20) => 
                           muxOutVector_4_20_port, A(19) => 
                           muxOutVector_4_19_port, A(18) => 
                           muxOutVector_4_18_port, A(17) => 
                           muxOutVector_4_17_port, A(16) => 
                           muxOutVector_4_16_port, A(15) => 
                           muxOutVector_4_15_port, A(14) => 
                           muxOutVector_4_14_port, A(13) => 
                           muxOutVector_4_13_port, A(12) => 
                           muxOutVector_4_12_port, A(11) => 
                           muxOutVector_4_11_port, A(10) => 
                           muxOutVector_4_10_port, A(9) => 
                           muxOutVector_4_9_port, A(8) => muxOutVector_4_8_port
                           , A(7) => muxOutVector_4_7_port, A(6) => 
                           muxOutVector_4_6_port, A(5) => muxOutVector_4_5_port
                           , A(4) => muxOutVector_4_4_port, A(3) => 
                           muxOutVector_4_3_port, A(2) => muxOutVector_4_2_port
                           , A(1) => muxOutVector_4_1_port, A(0) => 
                           muxOutVector_4_0_port, B(63) => sumVector_3_63_port,
                           B(62) => sumVector_3_62_port, B(61) => 
                           sumVector_3_61_port, B(60) => sumVector_3_60_port, 
                           B(59) => sumVector_3_59_port, B(58) => 
                           sumVector_3_58_port, B(57) => sumVector_3_57_port, 
                           B(56) => sumVector_3_56_port, B(55) => 
                           sumVector_3_55_port, B(54) => sumVector_3_54_port, 
                           B(53) => sumVector_3_53_port, B(52) => 
                           sumVector_3_52_port, B(51) => sumVector_3_51_port, 
                           B(50) => sumVector_3_50_port, B(49) => 
                           sumVector_3_49_port, B(48) => sumVector_3_48_port, 
                           B(47) => sumVector_3_47_port, B(46) => 
                           sumVector_3_46_port, B(45) => sumVector_3_45_port, 
                           B(44) => sumVector_3_44_port, B(43) => 
                           sumVector_3_43_port, B(42) => sumVector_3_42_port, 
                           B(41) => sumVector_3_41_port, B(40) => 
                           sumVector_3_40_port, B(39) => sumVector_3_39_port, 
                           B(38) => sumVector_3_38_port, B(37) => 
                           sumVector_3_37_port, B(36) => sumVector_3_36_port, 
                           B(35) => sumVector_3_35_port, B(34) => 
                           sumVector_3_34_port, B(33) => sumVector_3_33_port, 
                           B(32) => sumVector_3_32_port, B(31) => 
                           sumVector_3_31_port, B(30) => sumVector_3_30_port, 
                           B(29) => sumVector_3_29_port, B(28) => 
                           sumVector_3_28_port, B(27) => sumVector_3_27_port, 
                           B(26) => sumVector_3_26_port, B(25) => 
                           sumVector_3_25_port, B(24) => sumVector_3_24_port, 
                           B(23) => sumVector_3_23_port, B(22) => 
                           sumVector_3_22_port, B(21) => sumVector_3_21_port, 
                           B(20) => sumVector_3_20_port, B(19) => 
                           sumVector_3_19_port, B(18) => sumVector_3_18_port, 
                           B(17) => sumVector_3_17_port, B(16) => 
                           sumVector_3_16_port, B(15) => sumVector_3_15_port, 
                           B(14) => sumVector_3_14_port, B(13) => 
                           sumVector_3_13_port, B(12) => sumVector_3_12_port, 
                           B(11) => sumVector_3_11_port, B(10) => 
                           sumVector_3_10_port, B(9) => sumVector_3_9_port, 
                           B(8) => sumVector_3_8_port, B(7) => 
                           sumVector_3_7_port, B(6) => sumVector_3_6_port, B(5)
                           => sumVector_3_5_port, B(4) => sumVector_3_4_port, 
                           B(3) => sumVector_3_3_port, B(2) => 
                           sumVector_3_2_port, B(1) => sumVector_3_1_port, B(0)
                           => sumVector_3_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_4_63_port, S(62) => sumVector_4_62_port, 
                           S(61) => sumVector_4_61_port, S(60) => 
                           sumVector_4_60_port, S(59) => sumVector_4_59_port, 
                           S(58) => sumVector_4_58_port, S(57) => 
                           sumVector_4_57_port, S(56) => sumVector_4_56_port, 
                           S(55) => sumVector_4_55_port, S(54) => 
                           sumVector_4_54_port, S(53) => sumVector_4_53_port, 
                           S(52) => sumVector_4_52_port, S(51) => 
                           sumVector_4_51_port, S(50) => sumVector_4_50_port, 
                           S(49) => sumVector_4_49_port, S(48) => 
                           sumVector_4_48_port, S(47) => sumVector_4_47_port, 
                           S(46) => sumVector_4_46_port, S(45) => 
                           sumVector_4_45_port, S(44) => sumVector_4_44_port, 
                           S(43) => sumVector_4_43_port, S(42) => 
                           sumVector_4_42_port, S(41) => sumVector_4_41_port, 
                           S(40) => sumVector_4_40_port, S(39) => 
                           sumVector_4_39_port, S(38) => sumVector_4_38_port, 
                           S(37) => sumVector_4_37_port, S(36) => 
                           sumVector_4_36_port, S(35) => sumVector_4_35_port, 
                           S(34) => sumVector_4_34_port, S(33) => 
                           sumVector_4_33_port, S(32) => sumVector_4_32_port, 
                           S(31) => sumVector_4_31_port, S(30) => 
                           sumVector_4_30_port, S(29) => sumVector_4_29_port, 
                           S(28) => sumVector_4_28_port, S(27) => 
                           sumVector_4_27_port, S(26) => sumVector_4_26_port, 
                           S(25) => sumVector_4_25_port, S(24) => 
                           sumVector_4_24_port, S(23) => sumVector_4_23_port, 
                           S(22) => sumVector_4_22_port, S(21) => 
                           sumVector_4_21_port, S(20) => sumVector_4_20_port, 
                           S(19) => sumVector_4_19_port, S(18) => 
                           sumVector_4_18_port, S(17) => sumVector_4_17_port, 
                           S(16) => sumVector_4_16_port, S(15) => 
                           sumVector_4_15_port, S(14) => sumVector_4_14_port, 
                           S(13) => sumVector_4_13_port, S(12) => 
                           sumVector_4_12_port, S(11) => sumVector_4_11_port, 
                           S(10) => sumVector_4_10_port, S(9) => 
                           sumVector_4_9_port, S(8) => sumVector_4_8_port, S(7)
                           => sumVector_4_7_port, S(6) => sumVector_4_6_port, 
                           S(5) => sumVector_4_5_port, S(4) => 
                           sumVector_4_4_port, S(3) => sumVector_4_3_port, S(2)
                           => sumVector_4_2_port, S(1) => sumVector_4_1_port, 
                           S(0) => sumVector_4_0_port, Co => n_1039);
   mux_4 : MUX_5TO1_NBIT64_12 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n128, A1(62) => n129, 
                           A1(61) => n129, A1(60) => n127, A1(59) => n128, 
                           A1(58) => n129, A1(57) => n128, A1(56) => n129, 
                           A1(55) => n128, A1(54) => n129, A1(53) => n129, 
                           A1(52) => n128, A1(51) => n127, A1(50) => n128, 
                           A1(49) => n128, A1(48) => n128, A1(47) => n127, 
                           A1(46) => n128, A1(45) => n128, A1(44) => n127, 
                           A1(43) => n128, A1(42) => n127, A1(41) => n127, 
                           A1(40) => n127, A1(39) => n127, A1(38) => n379, 
                           A1(37) => n372, A1(36) => n365, A1(35) => n358, 
                           A1(34) => n351, A1(33) => n344, A1(32) => n337, 
                           A1(31) => n330, A1(30) => n323, A1(29) => n316, 
                           A1(28) => n309, A1(27) => n302, A1(26) => n295, 
                           A1(25) => n288, A1(24) => n281, A1(23) => n274, 
                           A1(22) => n267, A1(21) => n260, A1(20) => n253, 
                           A1(19) => n246, A1(18) => n239, A1(17) => n232, 
                           A1(16) => n225, A1(15) => n218, A1(14) => n211, 
                           A1(13) => n204, A1(12) => n197, A1(11) => n187, 
                           A1(10) => n181, A1(9) => n176, A1(8) => A(0), A1(7) 
                           => X_Logic0_port, A1(6) => X_Logic0_port, A1(5) => 
                           X_Logic0_port, A1(4) => X_Logic0_port, A1(3) => 
                           X_Logic0_port, A1(2) => X_Logic0_port, A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n529, A2(62) => n529, A2(61) => n529, A2(60) => n529
                           , A2(59) => n529, A2(58) => n529, A2(57) => n529, 
                           A2(56) => n529, A2(55) => n529, A2(54) => n529, 
                           A2(53) => n529, A2(52) => n529, A2(51) => n528, 
                           A2(50) => n528, A2(49) => n528, A2(48) => n528, 
                           A2(47) => n528, A2(46) => n528, A2(45) => n528, 
                           A2(44) => n528, A2(43) => n528, A2(42) => n528, 
                           A2(41) => n528, A2(40) => n528, A2(39) => n494, 
                           A2(38) => n490, A2(37) => n486, A2(36) => n482, 
                           A2(35) => n478, A2(34) => n474, A2(33) => n470, 
                           A2(32) => n466, A2(31) => n462, A2(30) => n458, 
                           A2(29) => n454, A2(28) => n450, A2(27) => n446, 
                           A2(26) => n442, A2(25) => n438, A2(24) => n434, 
                           A2(23) => n431, A2(22) => n427, A2(21) => n424, 
                           A2(20) => n421, A2(19) => n417, A2(18) => n413, 
                           A2(17) => n410, A2(16) => n406, A2(15) => n402, 
                           A2(14) => n105, A2(13) => n394, A2(12) => n392, 
                           A2(11) => n101, A2(10) => n387, A2(9) => n385, A2(8)
                           => n168, A2(7) => X_Logic0_port, A2(6) => 
                           X_Logic0_port, A2(5) => X_Logic0_port, A2(4) => 
                           X_Logic0_port, A2(3) => X_Logic0_port, A2(2) => 
                           X_Logic0_port, A2(1) => X_Logic0_port, A2(0) => 
                           X_Logic0_port, A3(63) => n162, A3(62) => n162, 
                           A3(61) => n162, A3(60) => n162, A3(59) => n162, 
                           A3(58) => n162, A3(57) => n557, A3(56) => n557, 
                           A3(55) => n557, A3(54) => n557, A3(53) => n557, 
                           A3(52) => n557, A3(51) => n557, A3(50) => n557, 
                           A3(49) => n557, A3(48) => n143, A3(47) => n143, 
                           A3(46) => n145, A3(45) => n144, A3(44) => n144, 
                           A3(43) => n145, A3(42) => n143, A3(41) => n144, 
                           A3(40) => n144, A3(39) => n375, A3(38) => n368, 
                           A3(37) => n361, A3(36) => n354, A3(35) => n347, 
                           A3(34) => n340, A3(33) => n333, A3(32) => n326, 
                           A3(31) => n319, A3(30) => n312, A3(29) => n305, 
                           A3(28) => n298, A3(27) => n291, A3(26) => n284, 
                           A3(25) => n277, A3(24) => n270, A3(23) => n263, 
                           A3(22) => n256, A3(21) => n249, A3(20) => n242, 
                           A3(19) => n235, A3(18) => n228, A3(17) => n221, 
                           A3(16) => n214, A3(15) => n207, A3(14) => n200, 
                           A3(13) => n193, A3(12) => n189, A3(11) => n180, 
                           A3(10) => n176, A3(9) => A(0), A3(8) => 
                           X_Logic0_port, A3(7) => X_Logic0_port, A3(6) => 
                           X_Logic0_port, A3(5) => X_Logic0_port, A3(4) => 
                           X_Logic0_port, A3(3) => X_Logic0_port, A3(2) => 
                           X_Logic0_port, A3(1) => X_Logic0_port, A3(0) => 
                           X_Logic0_port, A4(63) => n497, A4(62) => n497, 
                           A4(61) => n497, A4(60) => n497, A4(59) => n497, 
                           A4(58) => n497, A4(57) => n496, A4(56) => n496, 
                           A4(55) => n496, A4(54) => n496, A4(53) => n496, 
                           A4(52) => n496, A4(51) => n496, A4(50) => n496, 
                           A4(49) => n496, A4(48) => n496, A4(47) => n496, 
                           A4(46) => n503, A4(45) => n517, A4(44) => n515, 
                           A4(43) => n517, A4(42) => n516, A4(41) => n517, 
                           A4(40) => n492, A4(39) => n488, A4(38) => n484, 
                           A4(37) => n480, A4(36) => n476, A4(35) => n472, 
                           A4(34) => n468, A4(33) => n464, A4(32) => n460, 
                           A4(31) => n456, A4(30) => n452, A4(29) => n448, 
                           A4(28) => n444, A4(27) => n440, A4(26) => n436, 
                           A4(25) => n432, A4(24) => n429, A4(23) => n425, 
                           A4(22) => n422, A4(21) => n419, A4(20) => n415, 
                           A4(19) => n411, A4(18) => n408, A4(17) => n404, 
                           A4(16) => n400, A4(15) => n398, A4(14) => n396, 
                           A4(13) => n391, A4(12) => n388, A4(11) => n386, 
                           A4(10) => n99, A4(9) => n167, A4(8) => X_Logic0_port
                           , A4(7) => X_Logic0_port, A4(6) => X_Logic0_port, 
                           A4(5) => X_Logic0_port, A4(4) => X_Logic0_port, 
                           A4(3) => X_Logic0_port, A4(2) => X_Logic0_port, 
                           A4(1) => X_Logic0_port, A4(0) => X_Logic0_port, 
                           sel(2) => selVector_4_2_port, sel(1) => 
                           selVector_4_1_port, sel(0) => selVector_4_0_port, 
                           O(63) => muxOutVector_4_63_port, O(62) => 
                           muxOutVector_4_62_port, O(61) => 
                           muxOutVector_4_61_port, O(60) => 
                           muxOutVector_4_60_port, O(59) => 
                           muxOutVector_4_59_port, O(58) => 
                           muxOutVector_4_58_port, O(57) => 
                           muxOutVector_4_57_port, O(56) => 
                           muxOutVector_4_56_port, O(55) => 
                           muxOutVector_4_55_port, O(54) => 
                           muxOutVector_4_54_port, O(53) => 
                           muxOutVector_4_53_port, O(52) => 
                           muxOutVector_4_52_port, O(51) => 
                           muxOutVector_4_51_port, O(50) => 
                           muxOutVector_4_50_port, O(49) => 
                           muxOutVector_4_49_port, O(48) => 
                           muxOutVector_4_48_port, O(47) => 
                           muxOutVector_4_47_port, O(46) => 
                           muxOutVector_4_46_port, O(45) => 
                           muxOutVector_4_45_port, O(44) => 
                           muxOutVector_4_44_port, O(43) => 
                           muxOutVector_4_43_port, O(42) => 
                           muxOutVector_4_42_port, O(41) => 
                           muxOutVector_4_41_port, O(40) => 
                           muxOutVector_4_40_port, O(39) => 
                           muxOutVector_4_39_port, O(38) => 
                           muxOutVector_4_38_port, O(37) => 
                           muxOutVector_4_37_port, O(36) => 
                           muxOutVector_4_36_port, O(35) => 
                           muxOutVector_4_35_port, O(34) => 
                           muxOutVector_4_34_port, O(33) => 
                           muxOutVector_4_33_port, O(32) => 
                           muxOutVector_4_32_port, O(31) => 
                           muxOutVector_4_31_port, O(30) => 
                           muxOutVector_4_30_port, O(29) => 
                           muxOutVector_4_29_port, O(28) => 
                           muxOutVector_4_28_port, O(27) => 
                           muxOutVector_4_27_port, O(26) => 
                           muxOutVector_4_26_port, O(25) => 
                           muxOutVector_4_25_port, O(24) => 
                           muxOutVector_4_24_port, O(23) => 
                           muxOutVector_4_23_port, O(22) => 
                           muxOutVector_4_22_port, O(21) => 
                           muxOutVector_4_21_port, O(20) => 
                           muxOutVector_4_20_port, O(19) => 
                           muxOutVector_4_19_port, O(18) => 
                           muxOutVector_4_18_port, O(17) => 
                           muxOutVector_4_17_port, O(16) => 
                           muxOutVector_4_16_port, O(15) => 
                           muxOutVector_4_15_port, O(14) => 
                           muxOutVector_4_14_port, O(13) => 
                           muxOutVector_4_13_port, O(12) => 
                           muxOutVector_4_12_port, O(11) => 
                           muxOutVector_4_11_port, O(10) => 
                           muxOutVector_4_10_port, O(9) => 
                           muxOutVector_4_9_port, O(8) => muxOutVector_4_8_port
                           , O(7) => muxOutVector_4_7_port, O(6) => 
                           muxOutVector_4_6_port, O(5) => muxOutVector_4_5_port
                           , O(4) => muxOutVector_4_4_port, O(3) => 
                           muxOutVector_4_3_port, O(2) => muxOutVector_4_2_port
                           , O(1) => muxOutVector_4_1_port, O(0) => 
                           muxOutVector_4_0_port);
   eb_5 : BE_BLOCK_11 port map( b(2) => B(11), b(1) => B(10), b(0) => B(9), 
                           sel(2) => selVector_5_2_port, sel(1) => 
                           selVector_5_1_port, sel(0) => selVector_5_0_port);
   sum_5 : RCA_NBIT64_11 port map( A(63) => muxOutVector_5_63_port, A(62) => 
                           muxOutVector_5_62_port, A(61) => 
                           muxOutVector_5_61_port, A(60) => 
                           muxOutVector_5_60_port, A(59) => 
                           muxOutVector_5_59_port, A(58) => 
                           muxOutVector_5_58_port, A(57) => 
                           muxOutVector_5_57_port, A(56) => 
                           muxOutVector_5_56_port, A(55) => 
                           muxOutVector_5_55_port, A(54) => 
                           muxOutVector_5_54_port, A(53) => 
                           muxOutVector_5_53_port, A(52) => 
                           muxOutVector_5_52_port, A(51) => 
                           muxOutVector_5_51_port, A(50) => 
                           muxOutVector_5_50_port, A(49) => 
                           muxOutVector_5_49_port, A(48) => 
                           muxOutVector_5_48_port, A(47) => 
                           muxOutVector_5_47_port, A(46) => 
                           muxOutVector_5_46_port, A(45) => 
                           muxOutVector_5_45_port, A(44) => 
                           muxOutVector_5_44_port, A(43) => 
                           muxOutVector_5_43_port, A(42) => 
                           muxOutVector_5_42_port, A(41) => 
                           muxOutVector_5_41_port, A(40) => 
                           muxOutVector_5_40_port, A(39) => 
                           muxOutVector_5_39_port, A(38) => 
                           muxOutVector_5_38_port, A(37) => 
                           muxOutVector_5_37_port, A(36) => 
                           muxOutVector_5_36_port, A(35) => 
                           muxOutVector_5_35_port, A(34) => 
                           muxOutVector_5_34_port, A(33) => 
                           muxOutVector_5_33_port, A(32) => 
                           muxOutVector_5_32_port, A(31) => 
                           muxOutVector_5_31_port, A(30) => 
                           muxOutVector_5_30_port, A(29) => 
                           muxOutVector_5_29_port, A(28) => 
                           muxOutVector_5_28_port, A(27) => 
                           muxOutVector_5_27_port, A(26) => 
                           muxOutVector_5_26_port, A(25) => 
                           muxOutVector_5_25_port, A(24) => 
                           muxOutVector_5_24_port, A(23) => 
                           muxOutVector_5_23_port, A(22) => 
                           muxOutVector_5_22_port, A(21) => 
                           muxOutVector_5_21_port, A(20) => 
                           muxOutVector_5_20_port, A(19) => 
                           muxOutVector_5_19_port, A(18) => 
                           muxOutVector_5_18_port, A(17) => 
                           muxOutVector_5_17_port, A(16) => 
                           muxOutVector_5_16_port, A(15) => 
                           muxOutVector_5_15_port, A(14) => 
                           muxOutVector_5_14_port, A(13) => 
                           muxOutVector_5_13_port, A(12) => 
                           muxOutVector_5_12_port, A(11) => 
                           muxOutVector_5_11_port, A(10) => 
                           muxOutVector_5_10_port, A(9) => 
                           muxOutVector_5_9_port, A(8) => muxOutVector_5_8_port
                           , A(7) => muxOutVector_5_7_port, A(6) => 
                           muxOutVector_5_6_port, A(5) => muxOutVector_5_5_port
                           , A(4) => muxOutVector_5_4_port, A(3) => 
                           muxOutVector_5_3_port, A(2) => muxOutVector_5_2_port
                           , A(1) => muxOutVector_5_1_port, A(0) => 
                           muxOutVector_5_0_port, B(63) => sumVector_4_63_port,
                           B(62) => sumVector_4_62_port, B(61) => 
                           sumVector_4_61_port, B(60) => sumVector_4_60_port, 
                           B(59) => sumVector_4_59_port, B(58) => 
                           sumVector_4_58_port, B(57) => sumVector_4_57_port, 
                           B(56) => sumVector_4_56_port, B(55) => 
                           sumVector_4_55_port, B(54) => sumVector_4_54_port, 
                           B(53) => sumVector_4_53_port, B(52) => 
                           sumVector_4_52_port, B(51) => sumVector_4_51_port, 
                           B(50) => sumVector_4_50_port, B(49) => 
                           sumVector_4_49_port, B(48) => sumVector_4_48_port, 
                           B(47) => sumVector_4_47_port, B(46) => 
                           sumVector_4_46_port, B(45) => sumVector_4_45_port, 
                           B(44) => sumVector_4_44_port, B(43) => 
                           sumVector_4_43_port, B(42) => sumVector_4_42_port, 
                           B(41) => sumVector_4_41_port, B(40) => 
                           sumVector_4_40_port, B(39) => sumVector_4_39_port, 
                           B(38) => sumVector_4_38_port, B(37) => 
                           sumVector_4_37_port, B(36) => sumVector_4_36_port, 
                           B(35) => sumVector_4_35_port, B(34) => 
                           sumVector_4_34_port, B(33) => sumVector_4_33_port, 
                           B(32) => sumVector_4_32_port, B(31) => 
                           sumVector_4_31_port, B(30) => sumVector_4_30_port, 
                           B(29) => sumVector_4_29_port, B(28) => 
                           sumVector_4_28_port, B(27) => sumVector_4_27_port, 
                           B(26) => sumVector_4_26_port, B(25) => 
                           sumVector_4_25_port, B(24) => sumVector_4_24_port, 
                           B(23) => sumVector_4_23_port, B(22) => 
                           sumVector_4_22_port, B(21) => sumVector_4_21_port, 
                           B(20) => sumVector_4_20_port, B(19) => 
                           sumVector_4_19_port, B(18) => sumVector_4_18_port, 
                           B(17) => sumVector_4_17_port, B(16) => 
                           sumVector_4_16_port, B(15) => sumVector_4_15_port, 
                           B(14) => sumVector_4_14_port, B(13) => 
                           sumVector_4_13_port, B(12) => sumVector_4_12_port, 
                           B(11) => sumVector_4_11_port, B(10) => 
                           sumVector_4_10_port, B(9) => sumVector_4_9_port, 
                           B(8) => sumVector_4_8_port, B(7) => 
                           sumVector_4_7_port, B(6) => sumVector_4_6_port, B(5)
                           => sumVector_4_5_port, B(4) => sumVector_4_4_port, 
                           B(3) => sumVector_4_3_port, B(2) => 
                           sumVector_4_2_port, B(1) => sumVector_4_1_port, B(0)
                           => sumVector_4_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_5_63_port, S(62) => sumVector_5_62_port, 
                           S(61) => sumVector_5_61_port, S(60) => 
                           sumVector_5_60_port, S(59) => sumVector_5_59_port, 
                           S(58) => sumVector_5_58_port, S(57) => 
                           sumVector_5_57_port, S(56) => sumVector_5_56_port, 
                           S(55) => sumVector_5_55_port, S(54) => 
                           sumVector_5_54_port, S(53) => sumVector_5_53_port, 
                           S(52) => sumVector_5_52_port, S(51) => 
                           sumVector_5_51_port, S(50) => sumVector_5_50_port, 
                           S(49) => sumVector_5_49_port, S(48) => 
                           sumVector_5_48_port, S(47) => sumVector_5_47_port, 
                           S(46) => sumVector_5_46_port, S(45) => 
                           sumVector_5_45_port, S(44) => sumVector_5_44_port, 
                           S(43) => sumVector_5_43_port, S(42) => 
                           sumVector_5_42_port, S(41) => sumVector_5_41_port, 
                           S(40) => sumVector_5_40_port, S(39) => 
                           sumVector_5_39_port, S(38) => sumVector_5_38_port, 
                           S(37) => sumVector_5_37_port, S(36) => 
                           sumVector_5_36_port, S(35) => sumVector_5_35_port, 
                           S(34) => sumVector_5_34_port, S(33) => 
                           sumVector_5_33_port, S(32) => sumVector_5_32_port, 
                           S(31) => sumVector_5_31_port, S(30) => 
                           sumVector_5_30_port, S(29) => sumVector_5_29_port, 
                           S(28) => sumVector_5_28_port, S(27) => 
                           sumVector_5_27_port, S(26) => sumVector_5_26_port, 
                           S(25) => sumVector_5_25_port, S(24) => 
                           sumVector_5_24_port, S(23) => sumVector_5_23_port, 
                           S(22) => sumVector_5_22_port, S(21) => 
                           sumVector_5_21_port, S(20) => sumVector_5_20_port, 
                           S(19) => sumVector_5_19_port, S(18) => 
                           sumVector_5_18_port, S(17) => sumVector_5_17_port, 
                           S(16) => sumVector_5_16_port, S(15) => 
                           sumVector_5_15_port, S(14) => sumVector_5_14_port, 
                           S(13) => sumVector_5_13_port, S(12) => 
                           sumVector_5_12_port, S(11) => sumVector_5_11_port, 
                           S(10) => sumVector_5_10_port, S(9) => 
                           sumVector_5_9_port, S(8) => sumVector_5_8_port, S(7)
                           => sumVector_5_7_port, S(6) => sumVector_5_6_port, 
                           S(5) => sumVector_5_5_port, S(4) => 
                           sumVector_5_4_port, S(3) => sumVector_5_3_port, S(2)
                           => sumVector_5_2_port, S(1) => sumVector_5_1_port, 
                           S(0) => sumVector_5_0_port, Co => n_1040);
   mux_5 : MUX_5TO1_NBIT64_11 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n108, A1(62) => n108, 
                           A1(61) => n108, A1(60) => n108, A1(59) => n108, 
                           A1(58) => n108, A1(57) => n108, A1(56) => n108, 
                           A1(55) => n108, A1(54) => n108, A1(53) => n108, 
                           A1(52) => n107, A1(51) => n107, A1(50) => n107, 
                           A1(49) => n107, A1(48) => n107, A1(47) => n107, 
                           A1(46) => n107, A1(45) => n107, A1(44) => n107, 
                           A1(43) => n107, A1(42) => n107, A1(41) => n107, 
                           A1(40) => n375, A1(39) => n368, A1(38) => n361, 
                           A1(37) => n354, A1(36) => n347, A1(35) => n340, 
                           A1(34) => n333, A1(33) => n326, A1(32) => n319, 
                           A1(31) => n312, A1(30) => n305, A1(29) => n298, 
                           A1(28) => n291, A1(27) => n284, A1(26) => n277, 
                           A1(25) => n270, A1(24) => n263, A1(23) => n256, 
                           A1(22) => n249, A1(21) => n242, A1(20) => n235, 
                           A1(19) => n228, A1(18) => n221, A1(17) => n214, 
                           A1(16) => n207, A1(15) => n200, A1(14) => n193, 
                           A1(13) => n186, A1(12) => n179, A1(11) => n176, 
                           A1(10) => A(0), A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(63) => n532, A2(62) => n532, 
                           A2(61) => n532, A2(60) => n532, A2(59) => n532, 
                           A2(58) => n532, A2(57) => n532, A2(56) => n532, 
                           A2(55) => n532, A2(54) => n532, A2(53) => n532, 
                           A2(52) => n532, A2(51) => n531, A2(50) => n531, 
                           A2(49) => n531, A2(48) => n531, A2(47) => n531, 
                           A2(46) => n531, A2(45) => n531, A2(44) => n531, 
                           A2(43) => n531, A2(42) => n531, A2(41) => n494, 
                           A2(40) => n490, A2(39) => n486, A2(38) => n482, 
                           A2(37) => n478, A2(36) => n474, A2(35) => n470, 
                           A2(34) => n466, A2(33) => n462, A2(32) => n458, 
                           A2(31) => n454, A2(30) => n450, A2(29) => n446, 
                           A2(28) => n442, A2(27) => n438, A2(26) => n434, 
                           A2(25) => n431, A2(24) => n427, A2(23) => n424, 
                           A2(22) => n421, A2(21) => n417, A2(20) => n413, 
                           A2(19) => n410, A2(18) => n406, A2(17) => n402, 
                           A2(16) => n105, A2(15) => n394, A2(14) => n392, 
                           A2(13) => n389, A2(12) => n387, A2(11) => n383, 
                           A2(10) => n168, A2(9) => X_Logic0_port, A2(8) => 
                           X_Logic0_port, A2(7) => X_Logic0_port, A2(6) => 
                           X_Logic0_port, A2(5) => X_Logic0_port, A2(4) => 
                           X_Logic0_port, A2(3) => X_Logic0_port, A2(2) => 
                           X_Logic0_port, A2(1) => X_Logic0_port, A2(0) => 
                           X_Logic0_port, A3(63) => n160, A3(62) => n160, 
                           A3(61) => n160, A3(60) => n160, A3(59) => n160, 
                           A3(58) => n161, A3(57) => n161, A3(56) => n161, 
                           A3(55) => n161, A3(54) => n161, A3(53) => n161, 
                           A3(52) => n161, A3(51) => n161, A3(50) => n161, 
                           A3(49) => n161, A3(48) => n161, A3(47) => n161, 
                           A3(46) => n162, A3(45) => n162, A3(44) => n162, 
                           A3(43) => n162, A3(42) => n162, A3(41) => n376, 
                           A3(40) => n369, A3(39) => n362, A3(38) => n355, 
                           A3(37) => n348, A3(36) => n341, A3(35) => n334, 
                           A3(34) => n327, A3(33) => n320, A3(32) => n313, 
                           A3(31) => n306, A3(30) => n299, A3(29) => n292, 
                           A3(28) => n285, A3(27) => n278, A3(26) => n271, 
                           A3(25) => n264, A3(24) => n257, A3(23) => n250, 
                           A3(22) => n243, A3(21) => n236, A3(20) => n229, 
                           A3(19) => n222, A3(18) => n215, A3(17) => n208, 
                           A3(16) => n201, A3(15) => n194, A3(14) => n186, 
                           A3(13) => n182, A3(12) => n176, A3(11) => A(0), 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n499, A4(62) => 
                           n499, A4(61) => n499, A4(60) => n498, A4(59) => n498
                           , A4(58) => n498, A4(57) => n498, A4(56) => n498, 
                           A4(55) => n498, A4(54) => n498, A4(53) => n498, 
                           A4(52) => n498, A4(51) => n498, A4(50) => n498, 
                           A4(49) => n498, A4(48) => n497, A4(47) => n497, 
                           A4(46) => n497, A4(45) => n497, A4(44) => n497, 
                           A4(43) => n497, A4(42) => n492, A4(41) => n488, 
                           A4(40) => n484, A4(39) => n480, A4(38) => n476, 
                           A4(37) => n472, A4(36) => n468, A4(35) => n464, 
                           A4(34) => n460, A4(33) => n456, A4(32) => n452, 
                           A4(31) => n448, A4(30) => n444, A4(29) => n440, 
                           A4(28) => n436, A4(27) => n432, A4(26) => n429, 
                           A4(25) => n425, A4(24) => n422, A4(23) => n419, 
                           A4(22) => n415, A4(21) => n411, A4(20) => n408, 
                           A4(19) => n404, A4(18) => n400, A4(17) => n397, 
                           A4(16) => n394, A4(15) => n391, A4(14) => n100, 
                           A4(13) => n386, A4(12) => n385, A4(11) => n167, 
                           A4(10) => X_Logic0_port, A4(9) => X_Logic0_port, 
                           A4(8) => X_Logic0_port, A4(7) => X_Logic0_port, 
                           A4(6) => X_Logic0_port, A4(5) => X_Logic0_port, 
                           A4(4) => X_Logic0_port, A4(3) => X_Logic0_port, 
                           A4(2) => X_Logic0_port, A4(1) => X_Logic0_port, 
                           A4(0) => X_Logic0_port, sel(2) => selVector_5_2_port
                           , sel(1) => selVector_5_1_port, sel(0) => 
                           selVector_5_0_port, O(63) => muxOutVector_5_63_port,
                           O(62) => muxOutVector_5_62_port, O(61) => 
                           muxOutVector_5_61_port, O(60) => 
                           muxOutVector_5_60_port, O(59) => 
                           muxOutVector_5_59_port, O(58) => 
                           muxOutVector_5_58_port, O(57) => 
                           muxOutVector_5_57_port, O(56) => 
                           muxOutVector_5_56_port, O(55) => 
                           muxOutVector_5_55_port, O(54) => 
                           muxOutVector_5_54_port, O(53) => 
                           muxOutVector_5_53_port, O(52) => 
                           muxOutVector_5_52_port, O(51) => 
                           muxOutVector_5_51_port, O(50) => 
                           muxOutVector_5_50_port, O(49) => 
                           muxOutVector_5_49_port, O(48) => 
                           muxOutVector_5_48_port, O(47) => 
                           muxOutVector_5_47_port, O(46) => 
                           muxOutVector_5_46_port, O(45) => 
                           muxOutVector_5_45_port, O(44) => 
                           muxOutVector_5_44_port, O(43) => 
                           muxOutVector_5_43_port, O(42) => 
                           muxOutVector_5_42_port, O(41) => 
                           muxOutVector_5_41_port, O(40) => 
                           muxOutVector_5_40_port, O(39) => 
                           muxOutVector_5_39_port, O(38) => 
                           muxOutVector_5_38_port, O(37) => 
                           muxOutVector_5_37_port, O(36) => 
                           muxOutVector_5_36_port, O(35) => 
                           muxOutVector_5_35_port, O(34) => 
                           muxOutVector_5_34_port, O(33) => 
                           muxOutVector_5_33_port, O(32) => 
                           muxOutVector_5_32_port, O(31) => 
                           muxOutVector_5_31_port, O(30) => 
                           muxOutVector_5_30_port, O(29) => 
                           muxOutVector_5_29_port, O(28) => 
                           muxOutVector_5_28_port, O(27) => 
                           muxOutVector_5_27_port, O(26) => 
                           muxOutVector_5_26_port, O(25) => 
                           muxOutVector_5_25_port, O(24) => 
                           muxOutVector_5_24_port, O(23) => 
                           muxOutVector_5_23_port, O(22) => 
                           muxOutVector_5_22_port, O(21) => 
                           muxOutVector_5_21_port, O(20) => 
                           muxOutVector_5_20_port, O(19) => 
                           muxOutVector_5_19_port, O(18) => 
                           muxOutVector_5_18_port, O(17) => 
                           muxOutVector_5_17_port, O(16) => 
                           muxOutVector_5_16_port, O(15) => 
                           muxOutVector_5_15_port, O(14) => 
                           muxOutVector_5_14_port, O(13) => 
                           muxOutVector_5_13_port, O(12) => 
                           muxOutVector_5_12_port, O(11) => 
                           muxOutVector_5_11_port, O(10) => 
                           muxOutVector_5_10_port, O(9) => 
                           muxOutVector_5_9_port, O(8) => muxOutVector_5_8_port
                           , O(7) => muxOutVector_5_7_port, O(6) => 
                           muxOutVector_5_6_port, O(5) => muxOutVector_5_5_port
                           , O(4) => muxOutVector_5_4_port, O(3) => 
                           muxOutVector_5_3_port, O(2) => muxOutVector_5_2_port
                           , O(1) => muxOutVector_5_1_port, O(0) => 
                           muxOutVector_5_0_port);
   eb_6 : BE_BLOCK_10 port map( b(2) => B(13), b(1) => B(12), b(0) => B(11), 
                           sel(2) => selVector_6_2_port, sel(1) => 
                           selVector_6_1_port, sel(0) => selVector_6_0_port);
   sum_6 : RCA_NBIT64_10 port map( A(63) => muxOutVector_6_63_port, A(62) => 
                           muxOutVector_6_62_port, A(61) => 
                           muxOutVector_6_61_port, A(60) => 
                           muxOutVector_6_60_port, A(59) => 
                           muxOutVector_6_59_port, A(58) => 
                           muxOutVector_6_58_port, A(57) => 
                           muxOutVector_6_57_port, A(56) => 
                           muxOutVector_6_56_port, A(55) => 
                           muxOutVector_6_55_port, A(54) => 
                           muxOutVector_6_54_port, A(53) => 
                           muxOutVector_6_53_port, A(52) => 
                           muxOutVector_6_52_port, A(51) => 
                           muxOutVector_6_51_port, A(50) => 
                           muxOutVector_6_50_port, A(49) => 
                           muxOutVector_6_49_port, A(48) => 
                           muxOutVector_6_48_port, A(47) => 
                           muxOutVector_6_47_port, A(46) => 
                           muxOutVector_6_46_port, A(45) => 
                           muxOutVector_6_45_port, A(44) => 
                           muxOutVector_6_44_port, A(43) => 
                           muxOutVector_6_43_port, A(42) => 
                           muxOutVector_6_42_port, A(41) => 
                           muxOutVector_6_41_port, A(40) => 
                           muxOutVector_6_40_port, A(39) => 
                           muxOutVector_6_39_port, A(38) => 
                           muxOutVector_6_38_port, A(37) => 
                           muxOutVector_6_37_port, A(36) => 
                           muxOutVector_6_36_port, A(35) => 
                           muxOutVector_6_35_port, A(34) => 
                           muxOutVector_6_34_port, A(33) => 
                           muxOutVector_6_33_port, A(32) => 
                           muxOutVector_6_32_port, A(31) => 
                           muxOutVector_6_31_port, A(30) => 
                           muxOutVector_6_30_port, A(29) => 
                           muxOutVector_6_29_port, A(28) => 
                           muxOutVector_6_28_port, A(27) => 
                           muxOutVector_6_27_port, A(26) => 
                           muxOutVector_6_26_port, A(25) => 
                           muxOutVector_6_25_port, A(24) => 
                           muxOutVector_6_24_port, A(23) => 
                           muxOutVector_6_23_port, A(22) => 
                           muxOutVector_6_22_port, A(21) => 
                           muxOutVector_6_21_port, A(20) => 
                           muxOutVector_6_20_port, A(19) => 
                           muxOutVector_6_19_port, A(18) => 
                           muxOutVector_6_18_port, A(17) => 
                           muxOutVector_6_17_port, A(16) => 
                           muxOutVector_6_16_port, A(15) => 
                           muxOutVector_6_15_port, A(14) => 
                           muxOutVector_6_14_port, A(13) => 
                           muxOutVector_6_13_port, A(12) => 
                           muxOutVector_6_12_port, A(11) => 
                           muxOutVector_6_11_port, A(10) => 
                           muxOutVector_6_10_port, A(9) => 
                           muxOutVector_6_9_port, A(8) => muxOutVector_6_8_port
                           , A(7) => muxOutVector_6_7_port, A(6) => 
                           muxOutVector_6_6_port, A(5) => muxOutVector_6_5_port
                           , A(4) => muxOutVector_6_4_port, A(3) => 
                           muxOutVector_6_3_port, A(2) => muxOutVector_6_2_port
                           , A(1) => muxOutVector_6_1_port, A(0) => 
                           muxOutVector_6_0_port, B(63) => sumVector_5_63_port,
                           B(62) => sumVector_5_62_port, B(61) => 
                           sumVector_5_61_port, B(60) => sumVector_5_60_port, 
                           B(59) => sumVector_5_59_port, B(58) => 
                           sumVector_5_58_port, B(57) => sumVector_5_57_port, 
                           B(56) => sumVector_5_56_port, B(55) => 
                           sumVector_5_55_port, B(54) => sumVector_5_54_port, 
                           B(53) => sumVector_5_53_port, B(52) => 
                           sumVector_5_52_port, B(51) => sumVector_5_51_port, 
                           B(50) => sumVector_5_50_port, B(49) => 
                           sumVector_5_49_port, B(48) => sumVector_5_48_port, 
                           B(47) => sumVector_5_47_port, B(46) => 
                           sumVector_5_46_port, B(45) => sumVector_5_45_port, 
                           B(44) => sumVector_5_44_port, B(43) => 
                           sumVector_5_43_port, B(42) => sumVector_5_42_port, 
                           B(41) => sumVector_5_41_port, B(40) => 
                           sumVector_5_40_port, B(39) => sumVector_5_39_port, 
                           B(38) => sumVector_5_38_port, B(37) => 
                           sumVector_5_37_port, B(36) => sumVector_5_36_port, 
                           B(35) => sumVector_5_35_port, B(34) => 
                           sumVector_5_34_port, B(33) => sumVector_5_33_port, 
                           B(32) => sumVector_5_32_port, B(31) => 
                           sumVector_5_31_port, B(30) => sumVector_5_30_port, 
                           B(29) => sumVector_5_29_port, B(28) => 
                           sumVector_5_28_port, B(27) => sumVector_5_27_port, 
                           B(26) => sumVector_5_26_port, B(25) => 
                           sumVector_5_25_port, B(24) => sumVector_5_24_port, 
                           B(23) => sumVector_5_23_port, B(22) => 
                           sumVector_5_22_port, B(21) => sumVector_5_21_port, 
                           B(20) => sumVector_5_20_port, B(19) => 
                           sumVector_5_19_port, B(18) => sumVector_5_18_port, 
                           B(17) => sumVector_5_17_port, B(16) => 
                           sumVector_5_16_port, B(15) => sumVector_5_15_port, 
                           B(14) => sumVector_5_14_port, B(13) => 
                           sumVector_5_13_port, B(12) => sumVector_5_12_port, 
                           B(11) => sumVector_5_11_port, B(10) => 
                           sumVector_5_10_port, B(9) => sumVector_5_9_port, 
                           B(8) => sumVector_5_8_port, B(7) => 
                           sumVector_5_7_port, B(6) => sumVector_5_6_port, B(5)
                           => sumVector_5_5_port, B(4) => sumVector_5_4_port, 
                           B(3) => sumVector_5_3_port, B(2) => 
                           sumVector_5_2_port, B(1) => sumVector_5_1_port, B(0)
                           => sumVector_5_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_6_63_port, S(62) => sumVector_6_62_port, 
                           S(61) => sumVector_6_61_port, S(60) => 
                           sumVector_6_60_port, S(59) => sumVector_6_59_port, 
                           S(58) => sumVector_6_58_port, S(57) => 
                           sumVector_6_57_port, S(56) => sumVector_6_56_port, 
                           S(55) => sumVector_6_55_port, S(54) => 
                           sumVector_6_54_port, S(53) => sumVector_6_53_port, 
                           S(52) => sumVector_6_52_port, S(51) => 
                           sumVector_6_51_port, S(50) => sumVector_6_50_port, 
                           S(49) => sumVector_6_49_port, S(48) => 
                           sumVector_6_48_port, S(47) => sumVector_6_47_port, 
                           S(46) => sumVector_6_46_port, S(45) => 
                           sumVector_6_45_port, S(44) => sumVector_6_44_port, 
                           S(43) => sumVector_6_43_port, S(42) => 
                           sumVector_6_42_port, S(41) => sumVector_6_41_port, 
                           S(40) => sumVector_6_40_port, S(39) => 
                           sumVector_6_39_port, S(38) => sumVector_6_38_port, 
                           S(37) => sumVector_6_37_port, S(36) => 
                           sumVector_6_36_port, S(35) => sumVector_6_35_port, 
                           S(34) => sumVector_6_34_port, S(33) => 
                           sumVector_6_33_port, S(32) => sumVector_6_32_port, 
                           S(31) => sumVector_6_31_port, S(30) => 
                           sumVector_6_30_port, S(29) => sumVector_6_29_port, 
                           S(28) => sumVector_6_28_port, S(27) => 
                           sumVector_6_27_port, S(26) => sumVector_6_26_port, 
                           S(25) => sumVector_6_25_port, S(24) => 
                           sumVector_6_24_port, S(23) => sumVector_6_23_port, 
                           S(22) => sumVector_6_22_port, S(21) => 
                           sumVector_6_21_port, S(20) => sumVector_6_20_port, 
                           S(19) => sumVector_6_19_port, S(18) => 
                           sumVector_6_18_port, S(17) => sumVector_6_17_port, 
                           S(16) => sumVector_6_16_port, S(15) => 
                           sumVector_6_15_port, S(14) => sumVector_6_14_port, 
                           S(13) => sumVector_6_13_port, S(12) => 
                           sumVector_6_12_port, S(11) => sumVector_6_11_port, 
                           S(10) => sumVector_6_10_port, S(9) => 
                           sumVector_6_9_port, S(8) => sumVector_6_8_port, S(7)
                           => sumVector_6_7_port, S(6) => sumVector_6_6_port, 
                           S(5) => sumVector_6_5_port, S(4) => 
                           sumVector_6_4_port, S(3) => sumVector_6_3_port, S(2)
                           => sumVector_6_2_port, S(1) => sumVector_6_1_port, 
                           S(0) => sumVector_6_0_port, Co => n_1041);
   mux_6 : MUX_5TO1_NBIT64_10 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n110, A1(62) => n110, 
                           A1(61) => n110, A1(60) => n110, A1(59) => n110, 
                           A1(58) => n110, A1(57) => n110, A1(56) => n110, 
                           A1(55) => n110, A1(54) => n109, A1(53) => n109, 
                           A1(52) => n109, A1(51) => n109, A1(50) => n109, 
                           A1(49) => n109, A1(48) => n109, A1(47) => n109, 
                           A1(46) => n109, A1(45) => n109, A1(44) => n109, 
                           A1(43) => n108, A1(42) => n380, A1(41) => n373, 
                           A1(40) => n366, A1(39) => n359, A1(38) => n352, 
                           A1(37) => n345, A1(36) => n338, A1(35) => n331, 
                           A1(34) => n324, A1(33) => n317, A1(32) => n310, 
                           A1(31) => n303, A1(30) => n296, A1(29) => n289, 
                           A1(28) => n282, A1(27) => n275, A1(26) => n268, 
                           A1(25) => n261, A1(24) => n254, A1(23) => n247, 
                           A1(22) => n240, A1(21) => n233, A1(20) => n226, 
                           A1(19) => n219, A1(18) => n212, A1(17) => n205, 
                           A1(16) => n198, A1(15) => n186, A1(14) => n182, 
                           A1(13) => n176, A1(12) => A(0), A1(11) => 
                           X_Logic0_port, A1(10) => X_Logic0_port, A1(9) => 
                           X_Logic0_port, A1(8) => X_Logic0_port, A1(7) => 
                           X_Logic0_port, A1(6) => X_Logic0_port, A1(5) => 
                           X_Logic0_port, A1(4) => X_Logic0_port, A1(3) => 
                           X_Logic0_port, A1(2) => X_Logic0_port, A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n534, A2(62) => n534, A2(61) => n534, A2(60) => n534
                           , A2(59) => n534, A2(58) => n534, A2(57) => n534, 
                           A2(56) => n534, A2(55) => n534, A2(54) => n534, 
                           A2(53) => n533, A2(52) => n533, A2(51) => n533, 
                           A2(50) => n533, A2(49) => n533, A2(48) => n533, 
                           A2(47) => n533, A2(46) => n533, A2(45) => n533, 
                           A2(44) => n533, A2(43) => n494, A2(42) => n490, 
                           A2(41) => n486, A2(40) => n482, A2(39) => n478, 
                           A2(38) => n474, A2(37) => n470, A2(36) => n466, 
                           A2(35) => n462, A2(34) => n458, A2(33) => n454, 
                           A2(32) => n450, A2(31) => n446, A2(30) => n442, 
                           A2(29) => n438, A2(28) => n434, A2(27) => n431, 
                           A2(26) => n427, A2(25) => n424, A2(24) => n421, 
                           A2(23) => n417, A2(22) => n413, A2(21) => n410, 
                           A2(20) => n406, A2(19) => n402, A2(18) => n104, 
                           A2(17) => n394, A2(16) => n392, A2(15) => n101, 
                           A2(14) => n387, A2(13) => n99, A2(12) => n168, 
                           A2(11) => X_Logic0_port, A2(10) => X_Logic0_port, 
                           A2(9) => X_Logic0_port, A2(8) => X_Logic0_port, 
                           A2(7) => X_Logic0_port, A2(6) => X_Logic0_port, 
                           A2(5) => X_Logic0_port, A2(4) => X_Logic0_port, 
                           A2(3) => X_Logic0_port, A2(2) => X_Logic0_port, 
                           A2(1) => X_Logic0_port, A2(0) => X_Logic0_port, 
                           A3(63) => n158, A3(62) => n159, A3(61) => n159, 
                           A3(60) => n159, A3(59) => n159, A3(58) => n159, 
                           A3(57) => n159, A3(56) => n159, A3(55) => n159, 
                           A3(54) => n159, A3(53) => n159, A3(52) => n159, 
                           A3(51) => n159, A3(50) => n160, A3(49) => n160, 
                           A3(48) => n160, A3(47) => n160, A3(46) => n160, 
                           A3(45) => n160, A3(44) => n160, A3(43) => n380, 
                           A3(42) => n373, A3(41) => n366, A3(40) => n359, 
                           A3(39) => n352, A3(38) => n345, A3(37) => n338, 
                           A3(36) => n331, A3(35) => n324, A3(34) => n317, 
                           A3(33) => n310, A3(32) => n303, A3(31) => n296, 
                           A3(30) => n289, A3(29) => n282, A3(28) => n275, 
                           A3(27) => n268, A3(26) => n261, A3(25) => n254, 
                           A3(24) => n247, A3(23) => n240, A3(22) => n233, 
                           A3(21) => n226, A3(20) => n219, A3(19) => n212, 
                           A3(18) => n205, A3(17) => n198, A3(16) => n186, 
                           A3(15) => n182, A3(14) => n176, A3(13) => A(0), 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n500, A4(62) => 
                           n500, A4(61) => n500, A4(60) => n500, A4(59) => n500
                           , A4(58) => n500, A4(57) => n500, A4(56) => n500, 
                           A4(55) => n500, A4(54) => n500, A4(53) => n499, 
                           A4(52) => n499, A4(51) => n499, A4(50) => n499, 
                           A4(49) => n499, A4(48) => n499, A4(47) => n499, 
                           A4(46) => n499, A4(45) => n499, A4(44) => n492, 
                           A4(43) => n488, A4(42) => n484, A4(41) => n480, 
                           A4(40) => n476, A4(39) => n472, A4(38) => n468, 
                           A4(37) => n464, A4(36) => n460, A4(35) => n456, 
                           A4(34) => n452, A4(33) => n448, A4(32) => n444, 
                           A4(31) => n440, A4(30) => n436, A4(29) => n432, 
                           A4(28) => n429, A4(27) => n425, A4(26) => n422, 
                           A4(25) => n419, A4(24) => n415, A4(23) => n411, 
                           A4(22) => n408, A4(21) => n404, A4(20) => n400, 
                           A4(19) => n398, A4(18) => n396, A4(17) => n391, 
                           A4(16) => n388, A4(15) => n386, A4(14) => n99, 
                           A4(13) => n167, A4(12) => X_Logic0_port, A4(11) => 
                           X_Logic0_port, A4(10) => X_Logic0_port, A4(9) => 
                           X_Logic0_port, A4(8) => X_Logic0_port, A4(7) => 
                           X_Logic0_port, A4(6) => X_Logic0_port, A4(5) => 
                           X_Logic0_port, A4(4) => X_Logic0_port, A4(3) => 
                           X_Logic0_port, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_6_2_port, sel(1) => selVector_6_1_port, 
                           sel(0) => selVector_6_0_port, O(63) => 
                           muxOutVector_6_63_port, O(62) => 
                           muxOutVector_6_62_port, O(61) => 
                           muxOutVector_6_61_port, O(60) => 
                           muxOutVector_6_60_port, O(59) => 
                           muxOutVector_6_59_port, O(58) => 
                           muxOutVector_6_58_port, O(57) => 
                           muxOutVector_6_57_port, O(56) => 
                           muxOutVector_6_56_port, O(55) => 
                           muxOutVector_6_55_port, O(54) => 
                           muxOutVector_6_54_port, O(53) => 
                           muxOutVector_6_53_port, O(52) => 
                           muxOutVector_6_52_port, O(51) => 
                           muxOutVector_6_51_port, O(50) => 
                           muxOutVector_6_50_port, O(49) => 
                           muxOutVector_6_49_port, O(48) => 
                           muxOutVector_6_48_port, O(47) => 
                           muxOutVector_6_47_port, O(46) => 
                           muxOutVector_6_46_port, O(45) => 
                           muxOutVector_6_45_port, O(44) => 
                           muxOutVector_6_44_port, O(43) => 
                           muxOutVector_6_43_port, O(42) => 
                           muxOutVector_6_42_port, O(41) => 
                           muxOutVector_6_41_port, O(40) => 
                           muxOutVector_6_40_port, O(39) => 
                           muxOutVector_6_39_port, O(38) => 
                           muxOutVector_6_38_port, O(37) => 
                           muxOutVector_6_37_port, O(36) => 
                           muxOutVector_6_36_port, O(35) => 
                           muxOutVector_6_35_port, O(34) => 
                           muxOutVector_6_34_port, O(33) => 
                           muxOutVector_6_33_port, O(32) => 
                           muxOutVector_6_32_port, O(31) => 
                           muxOutVector_6_31_port, O(30) => 
                           muxOutVector_6_30_port, O(29) => 
                           muxOutVector_6_29_port, O(28) => 
                           muxOutVector_6_28_port, O(27) => 
                           muxOutVector_6_27_port, O(26) => 
                           muxOutVector_6_26_port, O(25) => 
                           muxOutVector_6_25_port, O(24) => 
                           muxOutVector_6_24_port, O(23) => 
                           muxOutVector_6_23_port, O(22) => 
                           muxOutVector_6_22_port, O(21) => 
                           muxOutVector_6_21_port, O(20) => 
                           muxOutVector_6_20_port, O(19) => 
                           muxOutVector_6_19_port, O(18) => 
                           muxOutVector_6_18_port, O(17) => 
                           muxOutVector_6_17_port, O(16) => 
                           muxOutVector_6_16_port, O(15) => 
                           muxOutVector_6_15_port, O(14) => 
                           muxOutVector_6_14_port, O(13) => 
                           muxOutVector_6_13_port, O(12) => 
                           muxOutVector_6_12_port, O(11) => 
                           muxOutVector_6_11_port, O(10) => 
                           muxOutVector_6_10_port, O(9) => 
                           muxOutVector_6_9_port, O(8) => muxOutVector_6_8_port
                           , O(7) => muxOutVector_6_7_port, O(6) => 
                           muxOutVector_6_6_port, O(5) => muxOutVector_6_5_port
                           , O(4) => muxOutVector_6_4_port, O(3) => 
                           muxOutVector_6_3_port, O(2) => muxOutVector_6_2_port
                           , O(1) => muxOutVector_6_1_port, O(0) => 
                           muxOutVector_6_0_port);
   eb_7 : BE_BLOCK_9 port map( b(2) => B(15), b(1) => B(14), b(0) => B(13), 
                           sel(2) => selVector_7_2_port, sel(1) => 
                           selVector_7_1_port, sel(0) => selVector_7_0_port);
   sum_7 : RCA_NBIT64_9 port map( A(63) => muxOutVector_7_63_port, A(62) => 
                           muxOutVector_7_62_port, A(61) => 
                           muxOutVector_7_61_port, A(60) => 
                           muxOutVector_7_60_port, A(59) => 
                           muxOutVector_7_59_port, A(58) => 
                           muxOutVector_7_58_port, A(57) => 
                           muxOutVector_7_57_port, A(56) => 
                           muxOutVector_7_56_port, A(55) => 
                           muxOutVector_7_55_port, A(54) => 
                           muxOutVector_7_54_port, A(53) => 
                           muxOutVector_7_53_port, A(52) => 
                           muxOutVector_7_52_port, A(51) => 
                           muxOutVector_7_51_port, A(50) => 
                           muxOutVector_7_50_port, A(49) => 
                           muxOutVector_7_49_port, A(48) => 
                           muxOutVector_7_48_port, A(47) => 
                           muxOutVector_7_47_port, A(46) => 
                           muxOutVector_7_46_port, A(45) => 
                           muxOutVector_7_45_port, A(44) => 
                           muxOutVector_7_44_port, A(43) => 
                           muxOutVector_7_43_port, A(42) => 
                           muxOutVector_7_42_port, A(41) => 
                           muxOutVector_7_41_port, A(40) => 
                           muxOutVector_7_40_port, A(39) => 
                           muxOutVector_7_39_port, A(38) => 
                           muxOutVector_7_38_port, A(37) => 
                           muxOutVector_7_37_port, A(36) => 
                           muxOutVector_7_36_port, A(35) => 
                           muxOutVector_7_35_port, A(34) => 
                           muxOutVector_7_34_port, A(33) => 
                           muxOutVector_7_33_port, A(32) => 
                           muxOutVector_7_32_port, A(31) => 
                           muxOutVector_7_31_port, A(30) => 
                           muxOutVector_7_30_port, A(29) => 
                           muxOutVector_7_29_port, A(28) => 
                           muxOutVector_7_28_port, A(27) => 
                           muxOutVector_7_27_port, A(26) => 
                           muxOutVector_7_26_port, A(25) => 
                           muxOutVector_7_25_port, A(24) => 
                           muxOutVector_7_24_port, A(23) => 
                           muxOutVector_7_23_port, A(22) => 
                           muxOutVector_7_22_port, A(21) => 
                           muxOutVector_7_21_port, A(20) => 
                           muxOutVector_7_20_port, A(19) => 
                           muxOutVector_7_19_port, A(18) => 
                           muxOutVector_7_18_port, A(17) => 
                           muxOutVector_7_17_port, A(16) => 
                           muxOutVector_7_16_port, A(15) => 
                           muxOutVector_7_15_port, A(14) => 
                           muxOutVector_7_14_port, A(13) => 
                           muxOutVector_7_13_port, A(12) => 
                           muxOutVector_7_12_port, A(11) => 
                           muxOutVector_7_11_port, A(10) => 
                           muxOutVector_7_10_port, A(9) => 
                           muxOutVector_7_9_port, A(8) => muxOutVector_7_8_port
                           , A(7) => muxOutVector_7_7_port, A(6) => 
                           muxOutVector_7_6_port, A(5) => muxOutVector_7_5_port
                           , A(4) => muxOutVector_7_4_port, A(3) => 
                           muxOutVector_7_3_port, A(2) => muxOutVector_7_2_port
                           , A(1) => muxOutVector_7_1_port, A(0) => 
                           muxOutVector_7_0_port, B(63) => sumVector_6_63_port,
                           B(62) => sumVector_6_62_port, B(61) => 
                           sumVector_6_61_port, B(60) => sumVector_6_60_port, 
                           B(59) => sumVector_6_59_port, B(58) => 
                           sumVector_6_58_port, B(57) => sumVector_6_57_port, 
                           B(56) => sumVector_6_56_port, B(55) => 
                           sumVector_6_55_port, B(54) => sumVector_6_54_port, 
                           B(53) => sumVector_6_53_port, B(52) => 
                           sumVector_6_52_port, B(51) => sumVector_6_51_port, 
                           B(50) => sumVector_6_50_port, B(49) => 
                           sumVector_6_49_port, B(48) => sumVector_6_48_port, 
                           B(47) => sumVector_6_47_port, B(46) => 
                           sumVector_6_46_port, B(45) => sumVector_6_45_port, 
                           B(44) => sumVector_6_44_port, B(43) => 
                           sumVector_6_43_port, B(42) => sumVector_6_42_port, 
                           B(41) => sumVector_6_41_port, B(40) => 
                           sumVector_6_40_port, B(39) => sumVector_6_39_port, 
                           B(38) => sumVector_6_38_port, B(37) => 
                           sumVector_6_37_port, B(36) => sumVector_6_36_port, 
                           B(35) => sumVector_6_35_port, B(34) => 
                           sumVector_6_34_port, B(33) => sumVector_6_33_port, 
                           B(32) => sumVector_6_32_port, B(31) => 
                           sumVector_6_31_port, B(30) => sumVector_6_30_port, 
                           B(29) => sumVector_6_29_port, B(28) => 
                           sumVector_6_28_port, B(27) => sumVector_6_27_port, 
                           B(26) => sumVector_6_26_port, B(25) => 
                           sumVector_6_25_port, B(24) => sumVector_6_24_port, 
                           B(23) => sumVector_6_23_port, B(22) => 
                           sumVector_6_22_port, B(21) => sumVector_6_21_port, 
                           B(20) => sumVector_6_20_port, B(19) => 
                           sumVector_6_19_port, B(18) => sumVector_6_18_port, 
                           B(17) => sumVector_6_17_port, B(16) => 
                           sumVector_6_16_port, B(15) => sumVector_6_15_port, 
                           B(14) => sumVector_6_14_port, B(13) => 
                           sumVector_6_13_port, B(12) => sumVector_6_12_port, 
                           B(11) => sumVector_6_11_port, B(10) => 
                           sumVector_6_10_port, B(9) => sumVector_6_9_port, 
                           B(8) => sumVector_6_8_port, B(7) => 
                           sumVector_6_7_port, B(6) => sumVector_6_6_port, B(5)
                           => sumVector_6_5_port, B(4) => sumVector_6_4_port, 
                           B(3) => sumVector_6_3_port, B(2) => 
                           sumVector_6_2_port, B(1) => sumVector_6_1_port, B(0)
                           => sumVector_6_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_7_63_port, S(62) => sumVector_7_62_port, 
                           S(61) => sumVector_7_61_port, S(60) => 
                           sumVector_7_60_port, S(59) => sumVector_7_59_port, 
                           S(58) => sumVector_7_58_port, S(57) => 
                           sumVector_7_57_port, S(56) => sumVector_7_56_port, 
                           S(55) => sumVector_7_55_port, S(54) => 
                           sumVector_7_54_port, S(53) => sumVector_7_53_port, 
                           S(52) => sumVector_7_52_port, S(51) => 
                           sumVector_7_51_port, S(50) => sumVector_7_50_port, 
                           S(49) => sumVector_7_49_port, S(48) => 
                           sumVector_7_48_port, S(47) => sumVector_7_47_port, 
                           S(46) => sumVector_7_46_port, S(45) => 
                           sumVector_7_45_port, S(44) => sumVector_7_44_port, 
                           S(43) => sumVector_7_43_port, S(42) => 
                           sumVector_7_42_port, S(41) => sumVector_7_41_port, 
                           S(40) => sumVector_7_40_port, S(39) => 
                           sumVector_7_39_port, S(38) => sumVector_7_38_port, 
                           S(37) => sumVector_7_37_port, S(36) => 
                           sumVector_7_36_port, S(35) => sumVector_7_35_port, 
                           S(34) => sumVector_7_34_port, S(33) => 
                           sumVector_7_33_port, S(32) => sumVector_7_32_port, 
                           S(31) => sumVector_7_31_port, S(30) => 
                           sumVector_7_30_port, S(29) => sumVector_7_29_port, 
                           S(28) => sumVector_7_28_port, S(27) => 
                           sumVector_7_27_port, S(26) => sumVector_7_26_port, 
                           S(25) => sumVector_7_25_port, S(24) => 
                           sumVector_7_24_port, S(23) => sumVector_7_23_port, 
                           S(22) => sumVector_7_22_port, S(21) => 
                           sumVector_7_21_port, S(20) => sumVector_7_20_port, 
                           S(19) => sumVector_7_19_port, S(18) => 
                           sumVector_7_18_port, S(17) => sumVector_7_17_port, 
                           S(16) => sumVector_7_16_port, S(15) => 
                           sumVector_7_15_port, S(14) => sumVector_7_14_port, 
                           S(13) => sumVector_7_13_port, S(12) => 
                           sumVector_7_12_port, S(11) => sumVector_7_11_port, 
                           S(10) => sumVector_7_10_port, S(9) => 
                           sumVector_7_9_port, S(8) => sumVector_7_8_port, S(7)
                           => sumVector_7_7_port, S(6) => sumVector_7_6_port, 
                           S(5) => sumVector_7_5_port, S(4) => 
                           sumVector_7_4_port, S(3) => sumVector_7_3_port, S(2)
                           => sumVector_7_2_port, S(1) => sumVector_7_1_port, 
                           S(0) => sumVector_7_0_port, Co => n_1042);
   mux_7 : MUX_5TO1_NBIT64_9 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n113, A1(62) => n113, 
                           A1(61) => n113, A1(60) => n112, A1(59) => n113, 
                           A1(58) => n113, A1(57) => n112, A1(56) => n112, 
                           A1(55) => n112, A1(54) => n112, A1(53) => n112, 
                           A1(52) => n112, A1(51) => n112, A1(50) => n112, 
                           A1(49) => n112, A1(48) => n111, A1(47) => n112, 
                           A1(46) => n112, A1(45) => n111, A1(44) => n379, 
                           A1(43) => n372, A1(42) => n365, A1(41) => n358, 
                           A1(40) => n351, A1(39) => n344, A1(38) => n337, 
                           A1(37) => n330, A1(36) => n323, A1(35) => n316, 
                           A1(34) => n309, A1(33) => n302, A1(32) => n295, 
                           A1(31) => n288, A1(30) => n281, A1(29) => n274, 
                           A1(28) => n267, A1(27) => n260, A1(26) => n253, 
                           A1(25) => n246, A1(24) => n239, A1(23) => n232, 
                           A1(22) => n225, A1(21) => n218, A1(20) => n211, 
                           A1(19) => n204, A1(18) => n197, A1(17) => n186, 
                           A1(16) => n182, A1(15) => n176, A1(14) => A(0), 
                           A1(13) => X_Logic0_port, A1(12) => X_Logic0_port, 
                           A1(11) => X_Logic0_port, A1(10) => X_Logic0_port, 
                           A1(9) => X_Logic0_port, A1(8) => X_Logic0_port, 
                           A1(7) => X_Logic0_port, A1(6) => X_Logic0_port, 
                           A1(5) => X_Logic0_port, A1(4) => X_Logic0_port, 
                           A1(3) => X_Logic0_port, A1(2) => X_Logic0_port, 
                           A1(1) => X_Logic0_port, A1(0) => X_Logic0_port, 
                           A2(63) => n537, A2(62) => n537, A2(61) => n537, 
                           A2(60) => n537, A2(59) => n537, A2(58) => n537, 
                           A2(57) => n537, A2(56) => n537, A2(55) => n537, 
                           A2(54) => n536, A2(53) => n536, A2(52) => n536, 
                           A2(51) => n536, A2(50) => n536, A2(49) => n536, 
                           A2(48) => n536, A2(47) => n536, A2(46) => n536, 
                           A2(45) => n494, A2(44) => n490, A2(43) => n486, 
                           A2(42) => n482, A2(41) => n478, A2(40) => n474, 
                           A2(39) => n470, A2(38) => n466, A2(37) => n462, 
                           A2(36) => n458, A2(35) => n454, A2(34) => n450, 
                           A2(33) => n446, A2(32) => n442, A2(31) => n438, 
                           A2(30) => n434, A2(29) => n431, A2(28) => n427, 
                           A2(27) => n424, A2(26) => n421, A2(25) => n417, 
                           A2(24) => n413, A2(23) => n410, A2(22) => n406, 
                           A2(21) => n402, A2(20) => n397, A2(19) => n396, 
                           A2(18) => n392, A2(17) => n389, A2(16) => n387, 
                           A2(15) => n383, A2(14) => n168, A2(13) => 
                           X_Logic0_port, A2(12) => X_Logic0_port, A2(11) => 
                           X_Logic0_port, A2(10) => X_Logic0_port, A2(9) => 
                           X_Logic0_port, A2(8) => X_Logic0_port, A2(7) => 
                           X_Logic0_port, A2(6) => X_Logic0_port, A2(5) => 
                           X_Logic0_port, A2(4) => X_Logic0_port, A2(3) => 
                           X_Logic0_port, A2(2) => X_Logic0_port, A2(1) => 
                           X_Logic0_port, A2(0) => X_Logic0_port, A3(63) => 
                           n157, A3(62) => n157, A3(61) => n157, A3(60) => n157
                           , A3(59) => n157, A3(58) => n157, A3(57) => n157, 
                           A3(56) => n158, A3(55) => n158, A3(54) => n158, 
                           A3(53) => n158, A3(52) => n158, A3(51) => n158, 
                           A3(50) => n158, A3(49) => n158, A3(48) => n158, 
                           A3(47) => n158, A3(46) => n158, A3(45) => n376, 
                           A3(44) => n369, A3(43) => n362, A3(42) => n355, 
                           A3(41) => n348, A3(40) => n341, A3(39) => n334, 
                           A3(38) => n327, A3(37) => n320, A3(36) => n313, 
                           A3(35) => n306, A3(34) => n299, A3(33) => n292, 
                           A3(32) => n285, A3(31) => n278, A3(30) => n271, 
                           A3(29) => n264, A3(28) => n257, A3(27) => n250, 
                           A3(26) => n243, A3(25) => n236, A3(24) => n229, 
                           A3(23) => n222, A3(22) => n215, A3(21) => n208, 
                           A3(20) => n201, A3(19) => n194, A3(18) => n186, 
                           A3(17) => n182, A3(16) => n176, A3(15) => A(0), 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n502, A4(62) => 
                           n502, A4(61) => n502, A4(60) => n501, A4(59) => n501
                           , A4(58) => n501, A4(57) => n501, A4(56) => n501, 
                           A4(55) => n501, A4(54) => n501, A4(53) => n501, 
                           A4(52) => n501, A4(51) => n501, A4(50) => n501, 
                           A4(49) => n501, A4(48) => n500, A4(47) => n500, 
                           A4(46) => n492, A4(45) => n488, A4(44) => n484, 
                           A4(43) => n480, A4(42) => n476, A4(41) => n472, 
                           A4(40) => n468, A4(39) => n464, A4(38) => n460, 
                           A4(37) => n456, A4(36) => n452, A4(35) => n448, 
                           A4(34) => n444, A4(33) => n440, A4(32) => n436, 
                           A4(31) => n432, A4(30) => n429, A4(29) => n425, 
                           A4(28) => n422, A4(27) => n419, A4(26) => n415, 
                           A4(25) => n411, A4(24) => n408, A4(23) => n404, 
                           A4(22) => n400, A4(21) => n104, A4(20) => n394, 
                           A4(19) => n391, A4(18) => n100, A4(17) => n386, 
                           A4(16) => n99, A4(15) => n167, A4(14) => 
                           X_Logic0_port, A4(13) => X_Logic0_port, A4(12) => 
                           X_Logic0_port, A4(11) => X_Logic0_port, A4(10) => 
                           X_Logic0_port, A4(9) => X_Logic0_port, A4(8) => 
                           X_Logic0_port, A4(7) => X_Logic0_port, A4(6) => 
                           X_Logic0_port, A4(5) => X_Logic0_port, A4(4) => 
                           X_Logic0_port, A4(3) => X_Logic0_port, A4(2) => 
                           X_Logic0_port, A4(1) => X_Logic0_port, A4(0) => 
                           X_Logic0_port, sel(2) => selVector_7_2_port, sel(1) 
                           => selVector_7_1_port, sel(0) => selVector_7_0_port,
                           O(63) => muxOutVector_7_63_port, O(62) => 
                           muxOutVector_7_62_port, O(61) => 
                           muxOutVector_7_61_port, O(60) => 
                           muxOutVector_7_60_port, O(59) => 
                           muxOutVector_7_59_port, O(58) => 
                           muxOutVector_7_58_port, O(57) => 
                           muxOutVector_7_57_port, O(56) => 
                           muxOutVector_7_56_port, O(55) => 
                           muxOutVector_7_55_port, O(54) => 
                           muxOutVector_7_54_port, O(53) => 
                           muxOutVector_7_53_port, O(52) => 
                           muxOutVector_7_52_port, O(51) => 
                           muxOutVector_7_51_port, O(50) => 
                           muxOutVector_7_50_port, O(49) => 
                           muxOutVector_7_49_port, O(48) => 
                           muxOutVector_7_48_port, O(47) => 
                           muxOutVector_7_47_port, O(46) => 
                           muxOutVector_7_46_port, O(45) => 
                           muxOutVector_7_45_port, O(44) => 
                           muxOutVector_7_44_port, O(43) => 
                           muxOutVector_7_43_port, O(42) => 
                           muxOutVector_7_42_port, O(41) => 
                           muxOutVector_7_41_port, O(40) => 
                           muxOutVector_7_40_port, O(39) => 
                           muxOutVector_7_39_port, O(38) => 
                           muxOutVector_7_38_port, O(37) => 
                           muxOutVector_7_37_port, O(36) => 
                           muxOutVector_7_36_port, O(35) => 
                           muxOutVector_7_35_port, O(34) => 
                           muxOutVector_7_34_port, O(33) => 
                           muxOutVector_7_33_port, O(32) => 
                           muxOutVector_7_32_port, O(31) => 
                           muxOutVector_7_31_port, O(30) => 
                           muxOutVector_7_30_port, O(29) => 
                           muxOutVector_7_29_port, O(28) => 
                           muxOutVector_7_28_port, O(27) => 
                           muxOutVector_7_27_port, O(26) => 
                           muxOutVector_7_26_port, O(25) => 
                           muxOutVector_7_25_port, O(24) => 
                           muxOutVector_7_24_port, O(23) => 
                           muxOutVector_7_23_port, O(22) => 
                           muxOutVector_7_22_port, O(21) => 
                           muxOutVector_7_21_port, O(20) => 
                           muxOutVector_7_20_port, O(19) => 
                           muxOutVector_7_19_port, O(18) => 
                           muxOutVector_7_18_port, O(17) => 
                           muxOutVector_7_17_port, O(16) => 
                           muxOutVector_7_16_port, O(15) => 
                           muxOutVector_7_15_port, O(14) => 
                           muxOutVector_7_14_port, O(13) => 
                           muxOutVector_7_13_port, O(12) => 
                           muxOutVector_7_12_port, O(11) => 
                           muxOutVector_7_11_port, O(10) => 
                           muxOutVector_7_10_port, O(9) => 
                           muxOutVector_7_9_port, O(8) => muxOutVector_7_8_port
                           , O(7) => muxOutVector_7_7_port, O(6) => 
                           muxOutVector_7_6_port, O(5) => muxOutVector_7_5_port
                           , O(4) => muxOutVector_7_4_port, O(3) => 
                           muxOutVector_7_3_port, O(2) => muxOutVector_7_2_port
                           , O(1) => muxOutVector_7_1_port, O(0) => 
                           muxOutVector_7_0_port);
   eb_8 : BE_BLOCK_8 port map( b(2) => B(17), b(1) => B(16), b(0) => B(15), 
                           sel(2) => selVector_8_2_port, sel(1) => 
                           selVector_8_1_port, sel(0) => selVector_8_0_port);
   sum_8 : RCA_NBIT64_8 port map( A(63) => muxOutVector_8_63_port, A(62) => 
                           muxOutVector_8_62_port, A(61) => 
                           muxOutVector_8_61_port, A(60) => 
                           muxOutVector_8_60_port, A(59) => 
                           muxOutVector_8_59_port, A(58) => 
                           muxOutVector_8_58_port, A(57) => 
                           muxOutVector_8_57_port, A(56) => 
                           muxOutVector_8_56_port, A(55) => 
                           muxOutVector_8_55_port, A(54) => 
                           muxOutVector_8_54_port, A(53) => 
                           muxOutVector_8_53_port, A(52) => 
                           muxOutVector_8_52_port, A(51) => 
                           muxOutVector_8_51_port, A(50) => 
                           muxOutVector_8_50_port, A(49) => 
                           muxOutVector_8_49_port, A(48) => 
                           muxOutVector_8_48_port, A(47) => 
                           muxOutVector_8_47_port, A(46) => 
                           muxOutVector_8_46_port, A(45) => 
                           muxOutVector_8_45_port, A(44) => 
                           muxOutVector_8_44_port, A(43) => 
                           muxOutVector_8_43_port, A(42) => 
                           muxOutVector_8_42_port, A(41) => 
                           muxOutVector_8_41_port, A(40) => 
                           muxOutVector_8_40_port, A(39) => 
                           muxOutVector_8_39_port, A(38) => 
                           muxOutVector_8_38_port, A(37) => 
                           muxOutVector_8_37_port, A(36) => 
                           muxOutVector_8_36_port, A(35) => 
                           muxOutVector_8_35_port, A(34) => 
                           muxOutVector_8_34_port, A(33) => 
                           muxOutVector_8_33_port, A(32) => 
                           muxOutVector_8_32_port, A(31) => 
                           muxOutVector_8_31_port, A(30) => 
                           muxOutVector_8_30_port, A(29) => 
                           muxOutVector_8_29_port, A(28) => 
                           muxOutVector_8_28_port, A(27) => 
                           muxOutVector_8_27_port, A(26) => 
                           muxOutVector_8_26_port, A(25) => 
                           muxOutVector_8_25_port, A(24) => 
                           muxOutVector_8_24_port, A(23) => 
                           muxOutVector_8_23_port, A(22) => 
                           muxOutVector_8_22_port, A(21) => 
                           muxOutVector_8_21_port, A(20) => 
                           muxOutVector_8_20_port, A(19) => 
                           muxOutVector_8_19_port, A(18) => 
                           muxOutVector_8_18_port, A(17) => 
                           muxOutVector_8_17_port, A(16) => 
                           muxOutVector_8_16_port, A(15) => 
                           muxOutVector_8_15_port, A(14) => 
                           muxOutVector_8_14_port, A(13) => 
                           muxOutVector_8_13_port, A(12) => 
                           muxOutVector_8_12_port, A(11) => 
                           muxOutVector_8_11_port, A(10) => 
                           muxOutVector_8_10_port, A(9) => 
                           muxOutVector_8_9_port, A(8) => muxOutVector_8_8_port
                           , A(7) => muxOutVector_8_7_port, A(6) => 
                           muxOutVector_8_6_port, A(5) => muxOutVector_8_5_port
                           , A(4) => muxOutVector_8_4_port, A(3) => 
                           muxOutVector_8_3_port, A(2) => muxOutVector_8_2_port
                           , A(1) => muxOutVector_8_1_port, A(0) => 
                           muxOutVector_8_0_port, B(63) => sumVector_7_63_port,
                           B(62) => sumVector_7_62_port, B(61) => 
                           sumVector_7_61_port, B(60) => sumVector_7_60_port, 
                           B(59) => sumVector_7_59_port, B(58) => 
                           sumVector_7_58_port, B(57) => sumVector_7_57_port, 
                           B(56) => sumVector_7_56_port, B(55) => 
                           sumVector_7_55_port, B(54) => sumVector_7_54_port, 
                           B(53) => sumVector_7_53_port, B(52) => 
                           sumVector_7_52_port, B(51) => sumVector_7_51_port, 
                           B(50) => sumVector_7_50_port, B(49) => 
                           sumVector_7_49_port, B(48) => sumVector_7_48_port, 
                           B(47) => sumVector_7_47_port, B(46) => 
                           sumVector_7_46_port, B(45) => sumVector_7_45_port, 
                           B(44) => sumVector_7_44_port, B(43) => 
                           sumVector_7_43_port, B(42) => sumVector_7_42_port, 
                           B(41) => sumVector_7_41_port, B(40) => 
                           sumVector_7_40_port, B(39) => sumVector_7_39_port, 
                           B(38) => sumVector_7_38_port, B(37) => 
                           sumVector_7_37_port, B(36) => sumVector_7_36_port, 
                           B(35) => sumVector_7_35_port, B(34) => 
                           sumVector_7_34_port, B(33) => sumVector_7_33_port, 
                           B(32) => sumVector_7_32_port, B(31) => 
                           sumVector_7_31_port, B(30) => sumVector_7_30_port, 
                           B(29) => sumVector_7_29_port, B(28) => 
                           sumVector_7_28_port, B(27) => sumVector_7_27_port, 
                           B(26) => sumVector_7_26_port, B(25) => 
                           sumVector_7_25_port, B(24) => sumVector_7_24_port, 
                           B(23) => sumVector_7_23_port, B(22) => 
                           sumVector_7_22_port, B(21) => sumVector_7_21_port, 
                           B(20) => sumVector_7_20_port, B(19) => 
                           sumVector_7_19_port, B(18) => sumVector_7_18_port, 
                           B(17) => sumVector_7_17_port, B(16) => 
                           sumVector_7_16_port, B(15) => sumVector_7_15_port, 
                           B(14) => sumVector_7_14_port, B(13) => 
                           sumVector_7_13_port, B(12) => sumVector_7_12_port, 
                           B(11) => sumVector_7_11_port, B(10) => 
                           sumVector_7_10_port, B(9) => sumVector_7_9_port, 
                           B(8) => sumVector_7_8_port, B(7) => 
                           sumVector_7_7_port, B(6) => sumVector_7_6_port, B(5)
                           => sumVector_7_5_port, B(4) => sumVector_7_4_port, 
                           B(3) => sumVector_7_3_port, B(2) => 
                           sumVector_7_2_port, B(1) => sumVector_7_1_port, B(0)
                           => sumVector_7_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_8_63_port, S(62) => sumVector_8_62_port, 
                           S(61) => sumVector_8_61_port, S(60) => 
                           sumVector_8_60_port, S(59) => sumVector_8_59_port, 
                           S(58) => sumVector_8_58_port, S(57) => 
                           sumVector_8_57_port, S(56) => sumVector_8_56_port, 
                           S(55) => sumVector_8_55_port, S(54) => 
                           sumVector_8_54_port, S(53) => sumVector_8_53_port, 
                           S(52) => sumVector_8_52_port, S(51) => 
                           sumVector_8_51_port, S(50) => sumVector_8_50_port, 
                           S(49) => sumVector_8_49_port, S(48) => 
                           sumVector_8_48_port, S(47) => sumVector_8_47_port, 
                           S(46) => sumVector_8_46_port, S(45) => 
                           sumVector_8_45_port, S(44) => sumVector_8_44_port, 
                           S(43) => sumVector_8_43_port, S(42) => 
                           sumVector_8_42_port, S(41) => sumVector_8_41_port, 
                           S(40) => sumVector_8_40_port, S(39) => 
                           sumVector_8_39_port, S(38) => sumVector_8_38_port, 
                           S(37) => sumVector_8_37_port, S(36) => 
                           sumVector_8_36_port, S(35) => sumVector_8_35_port, 
                           S(34) => sumVector_8_34_port, S(33) => 
                           sumVector_8_33_port, S(32) => sumVector_8_32_port, 
                           S(31) => sumVector_8_31_port, S(30) => 
                           sumVector_8_30_port, S(29) => sumVector_8_29_port, 
                           S(28) => sumVector_8_28_port, S(27) => 
                           sumVector_8_27_port, S(26) => sumVector_8_26_port, 
                           S(25) => sumVector_8_25_port, S(24) => 
                           sumVector_8_24_port, S(23) => sumVector_8_23_port, 
                           S(22) => sumVector_8_22_port, S(21) => 
                           sumVector_8_21_port, S(20) => sumVector_8_20_port, 
                           S(19) => sumVector_8_19_port, S(18) => 
                           sumVector_8_18_port, S(17) => sumVector_8_17_port, 
                           S(16) => sumVector_8_16_port, S(15) => 
                           sumVector_8_15_port, S(14) => sumVector_8_14_port, 
                           S(13) => sumVector_8_13_port, S(12) => 
                           sumVector_8_12_port, S(11) => sumVector_8_11_port, 
                           S(10) => sumVector_8_10_port, S(9) => 
                           sumVector_8_9_port, S(8) => sumVector_8_8_port, S(7)
                           => sumVector_8_7_port, S(6) => sumVector_8_6_port, 
                           S(5) => sumVector_8_5_port, S(4) => 
                           sumVector_8_4_port, S(3) => sumVector_8_3_port, S(2)
                           => sumVector_8_2_port, S(1) => sumVector_8_1_port, 
                           S(0) => sumVector_8_0_port, Co => n_1043);
   mux_8 : MUX_5TO1_NBIT64_8 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n115, A1(62) => n116, 
                           A1(61) => n116, A1(60) => n115, A1(59) => n115, 
                           A1(58) => n115, A1(57) => n115, A1(56) => n115, 
                           A1(55) => n115, A1(54) => n115, A1(53) => n115, 
                           A1(52) => n115, A1(51) => n114, A1(50) => n115, 
                           A1(49) => n115, A1(48) => n114, A1(47) => n114, 
                           A1(46) => n374, A1(45) => n367, A1(44) => n360, 
                           A1(43) => n353, A1(42) => n346, A1(41) => n339, 
                           A1(40) => n332, A1(39) => n325, A1(38) => n318, 
                           A1(37) => n311, A1(36) => n304, A1(35) => n297, 
                           A1(34) => n290, A1(33) => n283, A1(32) => n276, 
                           A1(31) => n269, A1(30) => n262, A1(29) => n255, 
                           A1(28) => n248, A1(27) => n241, A1(26) => n234, 
                           A1(25) => n227, A1(24) => n220, A1(23) => n213, 
                           A1(22) => n206, A1(21) => n199, A1(20) => n192, 
                           A1(19) => n186, A1(18) => n182, A1(17) => n176, 
                           A1(16) => A(0), A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(63) => n539, A2(62) => n539, 
                           A2(61) => n539, A2(60) => n539, A2(59) => n539, 
                           A2(58) => n539, A2(57) => n539, A2(56) => n539, 
                           A2(55) => n539, A2(54) => n539, A2(53) => n539, 
                           A2(52) => n538, A2(51) => n538, A2(50) => n538, 
                           A2(49) => n538, A2(48) => n538, A2(47) => n494, 
                           A2(46) => n490, A2(45) => n486, A2(44) => n482, 
                           A2(43) => n478, A2(42) => n474, A2(41) => n470, 
                           A2(40) => n466, A2(39) => n462, A2(38) => n458, 
                           A2(37) => n454, A2(36) => n450, A2(35) => n446, 
                           A2(34) => n442, A2(33) => n438, A2(32) => n434, 
                           A2(31) => n431, A2(30) => n427, A2(29) => n424, 
                           A2(28) => n421, A2(27) => n417, A2(26) => n413, 
                           A2(25) => n410, A2(24) => n405, A2(23) => n402, 
                           A2(22) => n105, A2(21) => n396, A2(20) => n392, 
                           A2(19) => n101, A2(18) => n387, A2(17) => n99, 
                           A2(16) => n168, A2(15) => X_Logic0_port, A2(14) => 
                           X_Logic0_port, A2(13) => X_Logic0_port, A2(12) => 
                           X_Logic0_port, A2(11) => X_Logic0_port, A2(10) => 
                           X_Logic0_port, A2(9) => X_Logic0_port, A2(8) => 
                           X_Logic0_port, A2(7) => X_Logic0_port, A2(6) => 
                           X_Logic0_port, A2(5) => X_Logic0_port, A2(4) => 
                           X_Logic0_port, A2(3) => X_Logic0_port, A2(2) => 
                           X_Logic0_port, A2(1) => X_Logic0_port, A2(0) => 
                           X_Logic0_port, A3(63) => n156, A3(62) => n156, 
                           A3(61) => n156, A3(60) => n156, A3(59) => n156, 
                           A3(58) => n156, A3(57) => n156, A3(56) => n156, 
                           A3(55) => n156, A3(54) => n156, A3(53) => n156, 
                           A3(52) => n157, A3(51) => n157, A3(50) => n157, 
                           A3(49) => n157, A3(48) => n157, A3(47) => n374, 
                           A3(46) => n367, A3(45) => n360, A3(44) => n353, 
                           A3(43) => n346, A3(42) => n339, A3(41) => n332, 
                           A3(40) => n325, A3(39) => n318, A3(38) => n311, 
                           A3(37) => n304, A3(36) => n297, A3(35) => n290, 
                           A3(34) => n283, A3(33) => n276, A3(32) => n269, 
                           A3(31) => n262, A3(30) => n255, A3(29) => n248, 
                           A3(28) => n241, A3(27) => n234, A3(26) => n227, 
                           A3(25) => n220, A3(24) => n213, A3(23) => n206, 
                           A3(22) => n199, A3(21) => n192, A3(20) => n186, 
                           A3(19) => n182, A3(18) => n176, A3(17) => A(0), 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n503, A4(62) => 
                           n503, A4(61) => n503, A4(60) => n503, A4(59) => n503
                           , A4(58) => n503, A4(57) => n502, A4(56) => n502, 
                           A4(55) => n502, A4(54) => n502, A4(53) => n502, 
                           A4(52) => n502, A4(51) => n502, A4(50) => n502, 
                           A4(49) => n502, A4(48) => n492, A4(47) => n488, 
                           A4(46) => n484, A4(45) => n480, A4(44) => n476, 
                           A4(43) => n472, A4(42) => n468, A4(41) => n464, 
                           A4(40) => n460, A4(39) => n456, A4(38) => n452, 
                           A4(37) => n448, A4(36) => n444, A4(35) => n440, 
                           A4(34) => n436, A4(33) => n432, A4(32) => n429, 
                           A4(31) => n425, A4(30) => n422, A4(29) => n419, 
                           A4(28) => n415, A4(27) => n411, A4(26) => n408, 
                           A4(25) => n404, A4(24) => n400, A4(23) => n397, 
                           A4(22) => n394, A4(21) => n391, A4(20) => n388, 
                           A4(19) => n386, A4(18) => n385, A4(17) => n167, 
                           A4(16) => X_Logic0_port, A4(15) => X_Logic0_port, 
                           A4(14) => X_Logic0_port, A4(13) => X_Logic0_port, 
                           A4(12) => X_Logic0_port, A4(11) => X_Logic0_port, 
                           A4(10) => X_Logic0_port, A4(9) => X_Logic0_port, 
                           A4(8) => X_Logic0_port, A4(7) => X_Logic0_port, 
                           A4(6) => X_Logic0_port, A4(5) => X_Logic0_port, 
                           A4(4) => X_Logic0_port, A4(3) => X_Logic0_port, 
                           A4(2) => X_Logic0_port, A4(1) => X_Logic0_port, 
                           A4(0) => X_Logic0_port, sel(2) => selVector_8_2_port
                           , sel(1) => selVector_8_1_port, sel(0) => 
                           selVector_8_0_port, O(63) => muxOutVector_8_63_port,
                           O(62) => muxOutVector_8_62_port, O(61) => 
                           muxOutVector_8_61_port, O(60) => 
                           muxOutVector_8_60_port, O(59) => 
                           muxOutVector_8_59_port, O(58) => 
                           muxOutVector_8_58_port, O(57) => 
                           muxOutVector_8_57_port, O(56) => 
                           muxOutVector_8_56_port, O(55) => 
                           muxOutVector_8_55_port, O(54) => 
                           muxOutVector_8_54_port, O(53) => 
                           muxOutVector_8_53_port, O(52) => 
                           muxOutVector_8_52_port, O(51) => 
                           muxOutVector_8_51_port, O(50) => 
                           muxOutVector_8_50_port, O(49) => 
                           muxOutVector_8_49_port, O(48) => 
                           muxOutVector_8_48_port, O(47) => 
                           muxOutVector_8_47_port, O(46) => 
                           muxOutVector_8_46_port, O(45) => 
                           muxOutVector_8_45_port, O(44) => 
                           muxOutVector_8_44_port, O(43) => 
                           muxOutVector_8_43_port, O(42) => 
                           muxOutVector_8_42_port, O(41) => 
                           muxOutVector_8_41_port, O(40) => 
                           muxOutVector_8_40_port, O(39) => 
                           muxOutVector_8_39_port, O(38) => 
                           muxOutVector_8_38_port, O(37) => 
                           muxOutVector_8_37_port, O(36) => 
                           muxOutVector_8_36_port, O(35) => 
                           muxOutVector_8_35_port, O(34) => 
                           muxOutVector_8_34_port, O(33) => 
                           muxOutVector_8_33_port, O(32) => 
                           muxOutVector_8_32_port, O(31) => 
                           muxOutVector_8_31_port, O(30) => 
                           muxOutVector_8_30_port, O(29) => 
                           muxOutVector_8_29_port, O(28) => 
                           muxOutVector_8_28_port, O(27) => 
                           muxOutVector_8_27_port, O(26) => 
                           muxOutVector_8_26_port, O(25) => 
                           muxOutVector_8_25_port, O(24) => 
                           muxOutVector_8_24_port, O(23) => 
                           muxOutVector_8_23_port, O(22) => 
                           muxOutVector_8_22_port, O(21) => 
                           muxOutVector_8_21_port, O(20) => 
                           muxOutVector_8_20_port, O(19) => 
                           muxOutVector_8_19_port, O(18) => 
                           muxOutVector_8_18_port, O(17) => 
                           muxOutVector_8_17_port, O(16) => 
                           muxOutVector_8_16_port, O(15) => 
                           muxOutVector_8_15_port, O(14) => 
                           muxOutVector_8_14_port, O(13) => 
                           muxOutVector_8_13_port, O(12) => 
                           muxOutVector_8_12_port, O(11) => 
                           muxOutVector_8_11_port, O(10) => 
                           muxOutVector_8_10_port, O(9) => 
                           muxOutVector_8_9_port, O(8) => muxOutVector_8_8_port
                           , O(7) => muxOutVector_8_7_port, O(6) => 
                           muxOutVector_8_6_port, O(5) => muxOutVector_8_5_port
                           , O(4) => muxOutVector_8_4_port, O(3) => 
                           muxOutVector_8_3_port, O(2) => muxOutVector_8_2_port
                           , O(1) => muxOutVector_8_1_port, O(0) => 
                           muxOutVector_8_0_port);
   eb_9 : BE_BLOCK_7 port map( b(2) => B(19), b(1) => B(18), b(0) => B(17), 
                           sel(2) => selVector_9_2_port, sel(1) => 
                           selVector_9_1_port, sel(0) => selVector_9_0_port);
   sum_9 : RCA_NBIT64_7 port map( A(63) => muxOutVector_9_63_port, A(62) => 
                           muxOutVector_9_62_port, A(61) => 
                           muxOutVector_9_61_port, A(60) => 
                           muxOutVector_9_60_port, A(59) => 
                           muxOutVector_9_59_port, A(58) => 
                           muxOutVector_9_58_port, A(57) => 
                           muxOutVector_9_57_port, A(56) => 
                           muxOutVector_9_56_port, A(55) => 
                           muxOutVector_9_55_port, A(54) => 
                           muxOutVector_9_54_port, A(53) => 
                           muxOutVector_9_53_port, A(52) => 
                           muxOutVector_9_52_port, A(51) => 
                           muxOutVector_9_51_port, A(50) => 
                           muxOutVector_9_50_port, A(49) => 
                           muxOutVector_9_49_port, A(48) => 
                           muxOutVector_9_48_port, A(47) => 
                           muxOutVector_9_47_port, A(46) => 
                           muxOutVector_9_46_port, A(45) => 
                           muxOutVector_9_45_port, A(44) => 
                           muxOutVector_9_44_port, A(43) => 
                           muxOutVector_9_43_port, A(42) => 
                           muxOutVector_9_42_port, A(41) => 
                           muxOutVector_9_41_port, A(40) => 
                           muxOutVector_9_40_port, A(39) => 
                           muxOutVector_9_39_port, A(38) => 
                           muxOutVector_9_38_port, A(37) => 
                           muxOutVector_9_37_port, A(36) => 
                           muxOutVector_9_36_port, A(35) => 
                           muxOutVector_9_35_port, A(34) => 
                           muxOutVector_9_34_port, A(33) => 
                           muxOutVector_9_33_port, A(32) => 
                           muxOutVector_9_32_port, A(31) => 
                           muxOutVector_9_31_port, A(30) => 
                           muxOutVector_9_30_port, A(29) => 
                           muxOutVector_9_29_port, A(28) => 
                           muxOutVector_9_28_port, A(27) => 
                           muxOutVector_9_27_port, A(26) => 
                           muxOutVector_9_26_port, A(25) => 
                           muxOutVector_9_25_port, A(24) => 
                           muxOutVector_9_24_port, A(23) => 
                           muxOutVector_9_23_port, A(22) => 
                           muxOutVector_9_22_port, A(21) => 
                           muxOutVector_9_21_port, A(20) => 
                           muxOutVector_9_20_port, A(19) => 
                           muxOutVector_9_19_port, A(18) => 
                           muxOutVector_9_18_port, A(17) => 
                           muxOutVector_9_17_port, A(16) => 
                           muxOutVector_9_16_port, A(15) => 
                           muxOutVector_9_15_port, A(14) => 
                           muxOutVector_9_14_port, A(13) => 
                           muxOutVector_9_13_port, A(12) => 
                           muxOutVector_9_12_port, A(11) => 
                           muxOutVector_9_11_port, A(10) => 
                           muxOutVector_9_10_port, A(9) => 
                           muxOutVector_9_9_port, A(8) => muxOutVector_9_8_port
                           , A(7) => muxOutVector_9_7_port, A(6) => 
                           muxOutVector_9_6_port, A(5) => muxOutVector_9_5_port
                           , A(4) => muxOutVector_9_4_port, A(3) => 
                           muxOutVector_9_3_port, A(2) => muxOutVector_9_2_port
                           , A(1) => muxOutVector_9_1_port, A(0) => 
                           muxOutVector_9_0_port, B(63) => sumVector_8_63_port,
                           B(62) => sumVector_8_62_port, B(61) => 
                           sumVector_8_61_port, B(60) => sumVector_8_60_port, 
                           B(59) => sumVector_8_59_port, B(58) => 
                           sumVector_8_58_port, B(57) => sumVector_8_57_port, 
                           B(56) => sumVector_8_56_port, B(55) => 
                           sumVector_8_55_port, B(54) => sumVector_8_54_port, 
                           B(53) => sumVector_8_53_port, B(52) => 
                           sumVector_8_52_port, B(51) => sumVector_8_51_port, 
                           B(50) => sumVector_8_50_port, B(49) => 
                           sumVector_8_49_port, B(48) => sumVector_8_48_port, 
                           B(47) => sumVector_8_47_port, B(46) => 
                           sumVector_8_46_port, B(45) => sumVector_8_45_port, 
                           B(44) => sumVector_8_44_port, B(43) => 
                           sumVector_8_43_port, B(42) => sumVector_8_42_port, 
                           B(41) => sumVector_8_41_port, B(40) => 
                           sumVector_8_40_port, B(39) => sumVector_8_39_port, 
                           B(38) => sumVector_8_38_port, B(37) => 
                           sumVector_8_37_port, B(36) => sumVector_8_36_port, 
                           B(35) => sumVector_8_35_port, B(34) => 
                           sumVector_8_34_port, B(33) => sumVector_8_33_port, 
                           B(32) => sumVector_8_32_port, B(31) => 
                           sumVector_8_31_port, B(30) => sumVector_8_30_port, 
                           B(29) => sumVector_8_29_port, B(28) => 
                           sumVector_8_28_port, B(27) => sumVector_8_27_port, 
                           B(26) => sumVector_8_26_port, B(25) => 
                           sumVector_8_25_port, B(24) => sumVector_8_24_port, 
                           B(23) => sumVector_8_23_port, B(22) => 
                           sumVector_8_22_port, B(21) => sumVector_8_21_port, 
                           B(20) => sumVector_8_20_port, B(19) => 
                           sumVector_8_19_port, B(18) => sumVector_8_18_port, 
                           B(17) => sumVector_8_17_port, B(16) => 
                           sumVector_8_16_port, B(15) => sumVector_8_15_port, 
                           B(14) => sumVector_8_14_port, B(13) => 
                           sumVector_8_13_port, B(12) => sumVector_8_12_port, 
                           B(11) => sumVector_8_11_port, B(10) => 
                           sumVector_8_10_port, B(9) => sumVector_8_9_port, 
                           B(8) => sumVector_8_8_port, B(7) => 
                           sumVector_8_7_port, B(6) => sumVector_8_6_port, B(5)
                           => sumVector_8_5_port, B(4) => sumVector_8_4_port, 
                           B(3) => sumVector_8_3_port, B(2) => 
                           sumVector_8_2_port, B(1) => sumVector_8_1_port, B(0)
                           => sumVector_8_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_9_63_port, S(62) => sumVector_9_62_port, 
                           S(61) => sumVector_9_61_port, S(60) => 
                           sumVector_9_60_port, S(59) => sumVector_9_59_port, 
                           S(58) => sumVector_9_58_port, S(57) => 
                           sumVector_9_57_port, S(56) => sumVector_9_56_port, 
                           S(55) => sumVector_9_55_port, S(54) => 
                           sumVector_9_54_port, S(53) => sumVector_9_53_port, 
                           S(52) => sumVector_9_52_port, S(51) => 
                           sumVector_9_51_port, S(50) => sumVector_9_50_port, 
                           S(49) => sumVector_9_49_port, S(48) => 
                           sumVector_9_48_port, S(47) => sumVector_9_47_port, 
                           S(46) => sumVector_9_46_port, S(45) => 
                           sumVector_9_45_port, S(44) => sumVector_9_44_port, 
                           S(43) => sumVector_9_43_port, S(42) => 
                           sumVector_9_42_port, S(41) => sumVector_9_41_port, 
                           S(40) => sumVector_9_40_port, S(39) => 
                           sumVector_9_39_port, S(38) => sumVector_9_38_port, 
                           S(37) => sumVector_9_37_port, S(36) => 
                           sumVector_9_36_port, S(35) => sumVector_9_35_port, 
                           S(34) => sumVector_9_34_port, S(33) => 
                           sumVector_9_33_port, S(32) => sumVector_9_32_port, 
                           S(31) => sumVector_9_31_port, S(30) => 
                           sumVector_9_30_port, S(29) => sumVector_9_29_port, 
                           S(28) => sumVector_9_28_port, S(27) => 
                           sumVector_9_27_port, S(26) => sumVector_9_26_port, 
                           S(25) => sumVector_9_25_port, S(24) => 
                           sumVector_9_24_port, S(23) => sumVector_9_23_port, 
                           S(22) => sumVector_9_22_port, S(21) => 
                           sumVector_9_21_port, S(20) => sumVector_9_20_port, 
                           S(19) => sumVector_9_19_port, S(18) => 
                           sumVector_9_18_port, S(17) => sumVector_9_17_port, 
                           S(16) => sumVector_9_16_port, S(15) => 
                           sumVector_9_15_port, S(14) => sumVector_9_14_port, 
                           S(13) => sumVector_9_13_port, S(12) => 
                           sumVector_9_12_port, S(11) => sumVector_9_11_port, 
                           S(10) => sumVector_9_10_port, S(9) => 
                           sumVector_9_9_port, S(8) => sumVector_9_8_port, S(7)
                           => sumVector_9_7_port, S(6) => sumVector_9_6_port, 
                           S(5) => sumVector_9_5_port, S(4) => 
                           sumVector_9_4_port, S(3) => sumVector_9_3_port, S(2)
                           => sumVector_9_2_port, S(1) => sumVector_9_1_port, 
                           S(0) => sumVector_9_0_port, Co => n_1044);
   mux_9 : MUX_5TO1_NBIT64_7 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n137, A1(62) => n137, 
                           A1(61) => n137, A1(60) => n136, A1(59) => n137, 
                           A1(58) => n137, A1(57) => n136, A1(56) => n136, 
                           A1(55) => n136, A1(54) => n136, A1(53) => n109, 
                           A1(52) => n116, A1(51) => n116, A1(50) => n116, 
                           A1(49) => n116, A1(48) => n380, A1(47) => n373, 
                           A1(46) => n366, A1(45) => n359, A1(44) => n352, 
                           A1(43) => n345, A1(42) => n338, A1(41) => n331, 
                           A1(40) => n324, A1(39) => n317, A1(38) => n310, 
                           A1(37) => n303, A1(36) => n296, A1(35) => n289, 
                           A1(34) => n282, A1(33) => n275, A1(32) => n268, 
                           A1(31) => n261, A1(30) => n254, A1(29) => n247, 
                           A1(28) => n240, A1(27) => n233, A1(26) => n226, 
                           A1(25) => n219, A1(24) => n212, A1(23) => n205, 
                           A1(22) => n198, A1(21) => n186, A1(20) => n182, 
                           A1(19) => n103, A1(18) => A(0), A1(17) => 
                           X_Logic0_port, A1(16) => X_Logic0_port, A1(15) => 
                           X_Logic0_port, A1(14) => X_Logic0_port, A1(13) => 
                           X_Logic0_port, A1(12) => X_Logic0_port, A1(11) => 
                           X_Logic0_port, A1(10) => X_Logic0_port, A1(9) => 
                           X_Logic0_port, A1(8) => X_Logic0_port, A1(7) => 
                           X_Logic0_port, A1(6) => X_Logic0_port, A1(5) => 
                           X_Logic0_port, A1(4) => X_Logic0_port, A1(3) => 
                           X_Logic0_port, A1(2) => X_Logic0_port, A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n517, A2(62) => n518, A2(61) => n517, A2(60) => n517
                           , A2(59) => n518, A2(58) => n518, A2(57) => n517, 
                           A2(56) => n518, A2(55) => n517, A2(54) => n517, 
                           A2(53) => n518, A2(52) => n517, A2(51) => n518, 
                           A2(50) => n539, A2(49) => n494, A2(48) => n490, 
                           A2(47) => n486, A2(46) => n482, A2(45) => n478, 
                           A2(44) => n474, A2(43) => n470, A2(42) => n466, 
                           A2(41) => n462, A2(40) => n458, A2(39) => n454, 
                           A2(38) => n450, A2(37) => n446, A2(36) => n442, 
                           A2(35) => n438, A2(34) => n434, A2(33) => n431, 
                           A2(32) => n427, A2(31) => n424, A2(30) => n421, 
                           A2(29) => n417, A2(28) => n413, A2(27) => n410, 
                           A2(26) => n405, A2(25) => n402, A2(24) => n104, 
                           A2(23) => n396, A2(22) => n392, A2(21) => n389, 
                           A2(20) => n387, A2(19) => n99, A2(18) => n168, 
                           A2(17) => X_Logic0_port, A2(16) => X_Logic0_port, 
                           A2(15) => X_Logic0_port, A2(14) => X_Logic0_port, 
                           A2(13) => X_Logic0_port, A2(12) => X_Logic0_port, 
                           A2(11) => X_Logic0_port, A2(10) => X_Logic0_port, 
                           A2(9) => X_Logic0_port, A2(8) => X_Logic0_port, 
                           A2(7) => X_Logic0_port, A2(6) => X_Logic0_port, 
                           A2(5) => X_Logic0_port, A2(4) => X_Logic0_port, 
                           A2(3) => X_Logic0_port, A2(2) => X_Logic0_port, 
                           A2(1) => X_Logic0_port, A2(0) => X_Logic0_port, 
                           A3(63) => n154, A3(62) => n154, A3(61) => n155, 
                           A3(60) => n155, A3(59) => n155, A3(58) => n155, 
                           A3(57) => n155, A3(56) => n155, A3(55) => n155, 
                           A3(54) => n155, A3(53) => n155, A3(52) => n155, 
                           A3(51) => n155, A3(50) => n155, A3(49) => n378, 
                           A3(48) => n371, A3(47) => n364, A3(46) => n357, 
                           A3(45) => n350, A3(44) => n343, A3(43) => n336, 
                           A3(42) => n329, A3(41) => n322, A3(40) => n315, 
                           A3(39) => n308, A3(38) => n301, A3(37) => n294, 
                           A3(36) => n287, A3(35) => n280, A3(34) => n273, 
                           A3(33) => n266, A3(32) => n259, A3(31) => n252, 
                           A3(30) => n245, A3(29) => n238, A3(28) => n231, 
                           A3(27) => n224, A3(26) => n217, A3(25) => n210, 
                           A3(24) => n203, A3(23) => n196, A3(22) => n186, 
                           A3(21) => n182, A3(20) => n176, A3(19) => A(0), 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n504, A4(62) => 
                           n504, A4(61) => n504, A4(60) => n504, A4(59) => n504
                           , A4(58) => n504, A4(57) => n504, A4(56) => n504, 
                           A4(55) => n503, A4(54) => n503, A4(53) => n503, 
                           A4(52) => n503, A4(51) => n503, A4(50) => n493, 
                           A4(49) => n489, A4(48) => n485, A4(47) => n481, 
                           A4(46) => n477, A4(45) => n473, A4(44) => n469, 
                           A4(43) => n465, A4(42) => n461, A4(41) => n457, 
                           A4(40) => n453, A4(39) => n449, A4(38) => n445, 
                           A4(37) => n441, A4(36) => n437, A4(35) => n433, 
                           A4(34) => n430, A4(33) => n426, A4(32) => n423, 
                           A4(31) => n420, A4(30) => n416, A4(29) => n412, 
                           A4(28) => n409, A4(27) => n404, A4(26) => n401, 
                           A4(25) => n398, A4(24) => n394, A4(23) => n391, 
                           A4(22) => n100, A4(21) => n386, A4(20) => n383, 
                           A4(19) => n167, A4(18) => X_Logic0_port, A4(17) => 
                           X_Logic0_port, A4(16) => X_Logic0_port, A4(15) => 
                           X_Logic0_port, A4(14) => X_Logic0_port, A4(13) => 
                           X_Logic0_port, A4(12) => X_Logic0_port, A4(11) => 
                           X_Logic0_port, A4(10) => X_Logic0_port, A4(9) => 
                           X_Logic0_port, A4(8) => X_Logic0_port, A4(7) => 
                           X_Logic0_port, A4(6) => X_Logic0_port, A4(5) => 
                           X_Logic0_port, A4(4) => X_Logic0_port, A4(3) => 
                           X_Logic0_port, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_9_2_port, sel(1) => selVector_9_1_port, 
                           sel(0) => selVector_9_0_port, O(63) => 
                           muxOutVector_9_63_port, O(62) => 
                           muxOutVector_9_62_port, O(61) => 
                           muxOutVector_9_61_port, O(60) => 
                           muxOutVector_9_60_port, O(59) => 
                           muxOutVector_9_59_port, O(58) => 
                           muxOutVector_9_58_port, O(57) => 
                           muxOutVector_9_57_port, O(56) => 
                           muxOutVector_9_56_port, O(55) => 
                           muxOutVector_9_55_port, O(54) => 
                           muxOutVector_9_54_port, O(53) => 
                           muxOutVector_9_53_port, O(52) => 
                           muxOutVector_9_52_port, O(51) => 
                           muxOutVector_9_51_port, O(50) => 
                           muxOutVector_9_50_port, O(49) => 
                           muxOutVector_9_49_port, O(48) => 
                           muxOutVector_9_48_port, O(47) => 
                           muxOutVector_9_47_port, O(46) => 
                           muxOutVector_9_46_port, O(45) => 
                           muxOutVector_9_45_port, O(44) => 
                           muxOutVector_9_44_port, O(43) => 
                           muxOutVector_9_43_port, O(42) => 
                           muxOutVector_9_42_port, O(41) => 
                           muxOutVector_9_41_port, O(40) => 
                           muxOutVector_9_40_port, O(39) => 
                           muxOutVector_9_39_port, O(38) => 
                           muxOutVector_9_38_port, O(37) => 
                           muxOutVector_9_37_port, O(36) => 
                           muxOutVector_9_36_port, O(35) => 
                           muxOutVector_9_35_port, O(34) => 
                           muxOutVector_9_34_port, O(33) => 
                           muxOutVector_9_33_port, O(32) => 
                           muxOutVector_9_32_port, O(31) => 
                           muxOutVector_9_31_port, O(30) => 
                           muxOutVector_9_30_port, O(29) => 
                           muxOutVector_9_29_port, O(28) => 
                           muxOutVector_9_28_port, O(27) => 
                           muxOutVector_9_27_port, O(26) => 
                           muxOutVector_9_26_port, O(25) => 
                           muxOutVector_9_25_port, O(24) => 
                           muxOutVector_9_24_port, O(23) => 
                           muxOutVector_9_23_port, O(22) => 
                           muxOutVector_9_22_port, O(21) => 
                           muxOutVector_9_21_port, O(20) => 
                           muxOutVector_9_20_port, O(19) => 
                           muxOutVector_9_19_port, O(18) => 
                           muxOutVector_9_18_port, O(17) => 
                           muxOutVector_9_17_port, O(16) => 
                           muxOutVector_9_16_port, O(15) => 
                           muxOutVector_9_15_port, O(14) => 
                           muxOutVector_9_14_port, O(13) => 
                           muxOutVector_9_13_port, O(12) => 
                           muxOutVector_9_12_port, O(11) => 
                           muxOutVector_9_11_port, O(10) => 
                           muxOutVector_9_10_port, O(9) => 
                           muxOutVector_9_9_port, O(8) => muxOutVector_9_8_port
                           , O(7) => muxOutVector_9_7_port, O(6) => 
                           muxOutVector_9_6_port, O(5) => muxOutVector_9_5_port
                           , O(4) => muxOutVector_9_4_port, O(3) => 
                           muxOutVector_9_3_port, O(2) => muxOutVector_9_2_port
                           , O(1) => muxOutVector_9_1_port, O(0) => 
                           muxOutVector_9_0_port);
   eb_10 : BE_BLOCK_6 port map( b(2) => B(21), b(1) => B(20), b(0) => B(19), 
                           sel(2) => selVector_10_2_port, sel(1) => 
                           selVector_10_1_port, sel(0) => selVector_10_0_port);
   sum_10 : RCA_NBIT64_6 port map( A(63) => muxOutVector_10_63_port, A(62) => 
                           muxOutVector_10_62_port, A(61) => 
                           muxOutVector_10_61_port, A(60) => 
                           muxOutVector_10_60_port, A(59) => 
                           muxOutVector_10_59_port, A(58) => 
                           muxOutVector_10_58_port, A(57) => 
                           muxOutVector_10_57_port, A(56) => 
                           muxOutVector_10_56_port, A(55) => 
                           muxOutVector_10_55_port, A(54) => 
                           muxOutVector_10_54_port, A(53) => 
                           muxOutVector_10_53_port, A(52) => 
                           muxOutVector_10_52_port, A(51) => 
                           muxOutVector_10_51_port, A(50) => 
                           muxOutVector_10_50_port, A(49) => 
                           muxOutVector_10_49_port, A(48) => 
                           muxOutVector_10_48_port, A(47) => 
                           muxOutVector_10_47_port, A(46) => 
                           muxOutVector_10_46_port, A(45) => 
                           muxOutVector_10_45_port, A(44) => 
                           muxOutVector_10_44_port, A(43) => 
                           muxOutVector_10_43_port, A(42) => 
                           muxOutVector_10_42_port, A(41) => 
                           muxOutVector_10_41_port, A(40) => 
                           muxOutVector_10_40_port, A(39) => 
                           muxOutVector_10_39_port, A(38) => 
                           muxOutVector_10_38_port, A(37) => 
                           muxOutVector_10_37_port, A(36) => 
                           muxOutVector_10_36_port, A(35) => 
                           muxOutVector_10_35_port, A(34) => 
                           muxOutVector_10_34_port, A(33) => 
                           muxOutVector_10_33_port, A(32) => 
                           muxOutVector_10_32_port, A(31) => 
                           muxOutVector_10_31_port, A(30) => 
                           muxOutVector_10_30_port, A(29) => 
                           muxOutVector_10_29_port, A(28) => 
                           muxOutVector_10_28_port, A(27) => 
                           muxOutVector_10_27_port, A(26) => 
                           muxOutVector_10_26_port, A(25) => 
                           muxOutVector_10_25_port, A(24) => 
                           muxOutVector_10_24_port, A(23) => 
                           muxOutVector_10_23_port, A(22) => 
                           muxOutVector_10_22_port, A(21) => 
                           muxOutVector_10_21_port, A(20) => 
                           muxOutVector_10_20_port, A(19) => 
                           muxOutVector_10_19_port, A(18) => 
                           muxOutVector_10_18_port, A(17) => 
                           muxOutVector_10_17_port, A(16) => 
                           muxOutVector_10_16_port, A(15) => 
                           muxOutVector_10_15_port, A(14) => 
                           muxOutVector_10_14_port, A(13) => 
                           muxOutVector_10_13_port, A(12) => 
                           muxOutVector_10_12_port, A(11) => 
                           muxOutVector_10_11_port, A(10) => 
                           muxOutVector_10_10_port, A(9) => 
                           muxOutVector_10_9_port, A(8) => 
                           muxOutVector_10_8_port, A(7) => 
                           muxOutVector_10_7_port, A(6) => 
                           muxOutVector_10_6_port, A(5) => 
                           muxOutVector_10_5_port, A(4) => 
                           muxOutVector_10_4_port, A(3) => 
                           muxOutVector_10_3_port, A(2) => 
                           muxOutVector_10_2_port, A(1) => 
                           muxOutVector_10_1_port, A(0) => 
                           muxOutVector_10_0_port, B(63) => sumVector_9_63_port
                           , B(62) => sumVector_9_62_port, B(61) => 
                           sumVector_9_61_port, B(60) => sumVector_9_60_port, 
                           B(59) => sumVector_9_59_port, B(58) => 
                           sumVector_9_58_port, B(57) => sumVector_9_57_port, 
                           B(56) => sumVector_9_56_port, B(55) => 
                           sumVector_9_55_port, B(54) => sumVector_9_54_port, 
                           B(53) => sumVector_9_53_port, B(52) => 
                           sumVector_9_52_port, B(51) => sumVector_9_51_port, 
                           B(50) => sumVector_9_50_port, B(49) => 
                           sumVector_9_49_port, B(48) => sumVector_9_48_port, 
                           B(47) => sumVector_9_47_port, B(46) => 
                           sumVector_9_46_port, B(45) => sumVector_9_45_port, 
                           B(44) => sumVector_9_44_port, B(43) => 
                           sumVector_9_43_port, B(42) => sumVector_9_42_port, 
                           B(41) => sumVector_9_41_port, B(40) => 
                           sumVector_9_40_port, B(39) => sumVector_9_39_port, 
                           B(38) => sumVector_9_38_port, B(37) => 
                           sumVector_9_37_port, B(36) => sumVector_9_36_port, 
                           B(35) => sumVector_9_35_port, B(34) => 
                           sumVector_9_34_port, B(33) => sumVector_9_33_port, 
                           B(32) => sumVector_9_32_port, B(31) => 
                           sumVector_9_31_port, B(30) => sumVector_9_30_port, 
                           B(29) => sumVector_9_29_port, B(28) => 
                           sumVector_9_28_port, B(27) => sumVector_9_27_port, 
                           B(26) => sumVector_9_26_port, B(25) => 
                           sumVector_9_25_port, B(24) => sumVector_9_24_port, 
                           B(23) => sumVector_9_23_port, B(22) => 
                           sumVector_9_22_port, B(21) => sumVector_9_21_port, 
                           B(20) => sumVector_9_20_port, B(19) => 
                           sumVector_9_19_port, B(18) => sumVector_9_18_port, 
                           B(17) => sumVector_9_17_port, B(16) => 
                           sumVector_9_16_port, B(15) => sumVector_9_15_port, 
                           B(14) => sumVector_9_14_port, B(13) => 
                           sumVector_9_13_port, B(12) => sumVector_9_12_port, 
                           B(11) => sumVector_9_11_port, B(10) => 
                           sumVector_9_10_port, B(9) => sumVector_9_9_port, 
                           B(8) => sumVector_9_8_port, B(7) => 
                           sumVector_9_7_port, B(6) => sumVector_9_6_port, B(5)
                           => sumVector_9_5_port, B(4) => sumVector_9_4_port, 
                           B(3) => sumVector_9_3_port, B(2) => 
                           sumVector_9_2_port, B(1) => sumVector_9_1_port, B(0)
                           => sumVector_9_0_port, Ci => X_Logic0_port, S(63) =>
                           sumVector_10_63_port, S(62) => sumVector_10_62_port,
                           S(61) => sumVector_10_61_port, S(60) => 
                           sumVector_10_60_port, S(59) => sumVector_10_59_port,
                           S(58) => sumVector_10_58_port, S(57) => 
                           sumVector_10_57_port, S(56) => sumVector_10_56_port,
                           S(55) => sumVector_10_55_port, S(54) => 
                           sumVector_10_54_port, S(53) => sumVector_10_53_port,
                           S(52) => sumVector_10_52_port, S(51) => 
                           sumVector_10_51_port, S(50) => sumVector_10_50_port,
                           S(49) => sumVector_10_49_port, S(48) => 
                           sumVector_10_48_port, S(47) => sumVector_10_47_port,
                           S(46) => sumVector_10_46_port, S(45) => 
                           sumVector_10_45_port, S(44) => sumVector_10_44_port,
                           S(43) => sumVector_10_43_port, S(42) => 
                           sumVector_10_42_port, S(41) => sumVector_10_41_port,
                           S(40) => sumVector_10_40_port, S(39) => 
                           sumVector_10_39_port, S(38) => sumVector_10_38_port,
                           S(37) => sumVector_10_37_port, S(36) => 
                           sumVector_10_36_port, S(35) => sumVector_10_35_port,
                           S(34) => sumVector_10_34_port, S(33) => 
                           sumVector_10_33_port, S(32) => sumVector_10_32_port,
                           S(31) => sumVector_10_31_port, S(30) => 
                           sumVector_10_30_port, S(29) => sumVector_10_29_port,
                           S(28) => sumVector_10_28_port, S(27) => 
                           sumVector_10_27_port, S(26) => sumVector_10_26_port,
                           S(25) => sumVector_10_25_port, S(24) => 
                           sumVector_10_24_port, S(23) => sumVector_10_23_port,
                           S(22) => sumVector_10_22_port, S(21) => 
                           sumVector_10_21_port, S(20) => sumVector_10_20_port,
                           S(19) => sumVector_10_19_port, S(18) => 
                           sumVector_10_18_port, S(17) => sumVector_10_17_port,
                           S(16) => sumVector_10_16_port, S(15) => 
                           sumVector_10_15_port, S(14) => sumVector_10_14_port,
                           S(13) => sumVector_10_13_port, S(12) => 
                           sumVector_10_12_port, S(11) => sumVector_10_11_port,
                           S(10) => sumVector_10_10_port, S(9) => 
                           sumVector_10_9_port, S(8) => sumVector_10_8_port, 
                           S(7) => sumVector_10_7_port, S(6) => 
                           sumVector_10_6_port, S(5) => sumVector_10_5_port, 
                           S(4) => sumVector_10_4_port, S(3) => 
                           sumVector_10_3_port, S(2) => sumVector_10_2_port, 
                           S(1) => sumVector_10_1_port, S(0) => 
                           sumVector_10_0_port, Co => n_1045);
   mux_10 : MUX_5TO1_NBIT64_6 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n121, A1(62) => n136, 
                           A1(61) => n121, A1(60) => n136, A1(59) => n136, 
                           A1(58) => n137, A1(57) => n136, A1(56) => n137, 
                           A1(55) => n136, A1(54) => n136, A1(53) => n137, 
                           A1(52) => n137, A1(51) => n136, A1(50) => n380, 
                           A1(49) => n373, A1(48) => n366, A1(47) => n359, 
                           A1(46) => n352, A1(45) => n345, A1(44) => n338, 
                           A1(43) => n331, A1(42) => n324, A1(41) => n317, 
                           A1(40) => n310, A1(39) => n303, A1(38) => n296, 
                           A1(37) => n289, A1(36) => n282, A1(35) => n275, 
                           A1(34) => n268, A1(33) => n261, A1(32) => n254, 
                           A1(31) => n247, A1(30) => n240, A1(29) => n233, 
                           A1(28) => n226, A1(27) => n219, A1(26) => n212, 
                           A1(25) => n205, A1(24) => n198, A1(23) => n186, 
                           A1(22) => n182, A1(21) => n103, A1(20) => A(0), 
                           A1(19) => X_Logic0_port, A1(18) => X_Logic0_port, 
                           A1(17) => X_Logic0_port, A1(16) => X_Logic0_port, 
                           A1(15) => X_Logic0_port, A1(14) => X_Logic0_port, 
                           A1(13) => X_Logic0_port, A1(12) => X_Logic0_port, 
                           A1(11) => X_Logic0_port, A1(10) => X_Logic0_port, 
                           A1(9) => X_Logic0_port, A1(8) => X_Logic0_port, 
                           A1(7) => X_Logic0_port, A1(6) => X_Logic0_port, 
                           A1(5) => X_Logic0_port, A1(4) => X_Logic0_port, 
                           A1(3) => X_Logic0_port, A1(2) => X_Logic0_port, 
                           A1(1) => X_Logic0_port, A1(0) => X_Logic0_port, 
                           A2(63) => n519, A2(62) => n519, A2(61) => n519, 
                           A2(60) => n521, A2(59) => n519, A2(58) => n519, 
                           A2(57) => n519, A2(56) => n518, A2(55) => n518, 
                           A2(54) => n518, A2(53) => n518, A2(52) => n517, 
                           A2(51) => n493, A2(50) => n489, A2(49) => n485, 
                           A2(48) => n481, A2(47) => n477, A2(46) => n473, 
                           A2(45) => n469, A2(44) => n465, A2(43) => n461, 
                           A2(42) => n457, A2(41) => n453, A2(40) => n449, 
                           A2(39) => n445, A2(38) => n441, A2(37) => n437, 
                           A2(36) => n433, A2(35) => n430, A2(34) => n426, 
                           A2(33) => n423, A2(32) => n420, A2(31) => n416, 
                           A2(30) => n412, A2(29) => n409, A2(28) => n405, 
                           A2(27) => n401, A2(26) => n105, A2(25) => n394, 
                           A2(24) => n392, A2(23) => n101, A2(22) => n387, 
                           A2(21) => n385, A2(20) => n168, A2(19) => 
                           X_Logic0_port, A2(18) => X_Logic0_port, A2(17) => 
                           X_Logic0_port, A2(16) => X_Logic0_port, A2(15) => 
                           X_Logic0_port, A2(14) => X_Logic0_port, A2(13) => 
                           X_Logic0_port, A2(12) => X_Logic0_port, A2(11) => 
                           X_Logic0_port, A2(10) => X_Logic0_port, A2(9) => 
                           X_Logic0_port, A2(8) => X_Logic0_port, A2(7) => 
                           X_Logic0_port, A2(6) => X_Logic0_port, A2(5) => 
                           X_Logic0_port, A2(4) => X_Logic0_port, A2(3) => 
                           X_Logic0_port, A2(2) => X_Logic0_port, A2(1) => 
                           X_Logic0_port, A2(0) => X_Logic0_port, A3(63) => 
                           n153, A3(62) => n153, A3(61) => n154, A3(60) => n154
                           , A3(59) => n154, A3(58) => n154, A3(57) => n154, 
                           A3(56) => n154, A3(55) => n154, A3(54) => n154, 
                           A3(53) => n154, A3(52) => n154, A3(51) => n377, 
                           A3(50) => n370, A3(49) => n363, A3(48) => n356, 
                           A3(47) => n349, A3(46) => n342, A3(45) => n335, 
                           A3(44) => n328, A3(43) => n321, A3(42) => n314, 
                           A3(41) => n307, A3(40) => n300, A3(39) => n293, 
                           A3(38) => n286, A3(37) => n279, A3(36) => n272, 
                           A3(35) => n265, A3(34) => n258, A3(33) => n251, 
                           A3(32) => n244, A3(31) => n237, A3(30) => n230, 
                           A3(29) => n223, A3(28) => n216, A3(27) => n209, 
                           A3(26) => n202, A3(25) => n195, A3(24) => n186, 
                           A3(23) => n182, A3(22) => n176, A3(21) => A(0), 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n505, A4(62) => 
                           n505, A4(61) => n505, A4(60) => n505, A4(59) => n505
                           , A4(58) => n505, A4(57) => n505, A4(56) => n504, 
                           A4(55) => n504, A4(54) => n504, A4(53) => n504, 
                           A4(52) => n493, A4(51) => n489, A4(50) => n485, 
                           A4(49) => n481, A4(48) => n477, A4(47) => n473, 
                           A4(46) => n469, A4(45) => n465, A4(44) => n461, 
                           A4(43) => n457, A4(42) => n453, A4(41) => n449, 
                           A4(40) => n445, A4(39) => n441, A4(38) => n437, 
                           A4(37) => n433, A4(36) => n430, A4(35) => n426, 
                           A4(34) => n423, A4(33) => n420, A4(32) => n416, 
                           A4(31) => n412, A4(30) => n409, A4(29) => n405, 
                           A4(28) => n401, A4(27) => n397, A4(26) => n396, 
                           A4(25) => n392, A4(24) => n388, A4(23) => n387, 
                           A4(22) => n99, A4(21) => n167, A4(20) => 
                           X_Logic0_port, A4(19) => X_Logic0_port, A4(18) => 
                           X_Logic0_port, A4(17) => X_Logic0_port, A4(16) => 
                           X_Logic0_port, A4(15) => X_Logic0_port, A4(14) => 
                           X_Logic0_port, A4(13) => X_Logic0_port, A4(12) => 
                           X_Logic0_port, A4(11) => X_Logic0_port, A4(10) => 
                           X_Logic0_port, A4(9) => X_Logic0_port, A4(8) => 
                           X_Logic0_port, A4(7) => X_Logic0_port, A4(6) => 
                           X_Logic0_port, A4(5) => X_Logic0_port, A4(4) => 
                           X_Logic0_port, A4(3) => X_Logic0_port, A4(2) => 
                           X_Logic0_port, A4(1) => X_Logic0_port, A4(0) => 
                           X_Logic0_port, sel(2) => selVector_10_2_port, sel(1)
                           => selVector_10_1_port, sel(0) => 
                           selVector_10_0_port, O(63) => 
                           muxOutVector_10_63_port, O(62) => 
                           muxOutVector_10_62_port, O(61) => 
                           muxOutVector_10_61_port, O(60) => 
                           muxOutVector_10_60_port, O(59) => 
                           muxOutVector_10_59_port, O(58) => 
                           muxOutVector_10_58_port, O(57) => 
                           muxOutVector_10_57_port, O(56) => 
                           muxOutVector_10_56_port, O(55) => 
                           muxOutVector_10_55_port, O(54) => 
                           muxOutVector_10_54_port, O(53) => 
                           muxOutVector_10_53_port, O(52) => 
                           muxOutVector_10_52_port, O(51) => 
                           muxOutVector_10_51_port, O(50) => 
                           muxOutVector_10_50_port, O(49) => 
                           muxOutVector_10_49_port, O(48) => 
                           muxOutVector_10_48_port, O(47) => 
                           muxOutVector_10_47_port, O(46) => 
                           muxOutVector_10_46_port, O(45) => 
                           muxOutVector_10_45_port, O(44) => 
                           muxOutVector_10_44_port, O(43) => 
                           muxOutVector_10_43_port, O(42) => 
                           muxOutVector_10_42_port, O(41) => 
                           muxOutVector_10_41_port, O(40) => 
                           muxOutVector_10_40_port, O(39) => 
                           muxOutVector_10_39_port, O(38) => 
                           muxOutVector_10_38_port, O(37) => 
                           muxOutVector_10_37_port, O(36) => 
                           muxOutVector_10_36_port, O(35) => 
                           muxOutVector_10_35_port, O(34) => 
                           muxOutVector_10_34_port, O(33) => 
                           muxOutVector_10_33_port, O(32) => 
                           muxOutVector_10_32_port, O(31) => 
                           muxOutVector_10_31_port, O(30) => 
                           muxOutVector_10_30_port, O(29) => 
                           muxOutVector_10_29_port, O(28) => 
                           muxOutVector_10_28_port, O(27) => 
                           muxOutVector_10_27_port, O(26) => 
                           muxOutVector_10_26_port, O(25) => 
                           muxOutVector_10_25_port, O(24) => 
                           muxOutVector_10_24_port, O(23) => 
                           muxOutVector_10_23_port, O(22) => 
                           muxOutVector_10_22_port, O(21) => 
                           muxOutVector_10_21_port, O(20) => 
                           muxOutVector_10_20_port, O(19) => 
                           muxOutVector_10_19_port, O(18) => 
                           muxOutVector_10_18_port, O(17) => 
                           muxOutVector_10_17_port, O(16) => 
                           muxOutVector_10_16_port, O(15) => 
                           muxOutVector_10_15_port, O(14) => 
                           muxOutVector_10_14_port, O(13) => 
                           muxOutVector_10_13_port, O(12) => 
                           muxOutVector_10_12_port, O(11) => 
                           muxOutVector_10_11_port, O(10) => 
                           muxOutVector_10_10_port, O(9) => 
                           muxOutVector_10_9_port, O(8) => 
                           muxOutVector_10_8_port, O(7) => 
                           muxOutVector_10_7_port, O(6) => 
                           muxOutVector_10_6_port, O(5) => 
                           muxOutVector_10_5_port, O(4) => 
                           muxOutVector_10_4_port, O(3) => 
                           muxOutVector_10_3_port, O(2) => 
                           muxOutVector_10_2_port, O(1) => 
                           muxOutVector_10_1_port, O(0) => 
                           muxOutVector_10_0_port);
   eb_11 : BE_BLOCK_5 port map( b(2) => B(23), b(1) => B(22), b(0) => B(21), 
                           sel(2) => selVector_11_2_port, sel(1) => 
                           selVector_11_1_port, sel(0) => selVector_11_0_port);
   sum_11 : RCA_NBIT64_5 port map( A(63) => muxOutVector_11_63_port, A(62) => 
                           muxOutVector_11_62_port, A(61) => 
                           muxOutVector_11_61_port, A(60) => 
                           muxOutVector_11_60_port, A(59) => 
                           muxOutVector_11_59_port, A(58) => 
                           muxOutVector_11_58_port, A(57) => 
                           muxOutVector_11_57_port, A(56) => 
                           muxOutVector_11_56_port, A(55) => 
                           muxOutVector_11_55_port, A(54) => 
                           muxOutVector_11_54_port, A(53) => 
                           muxOutVector_11_53_port, A(52) => 
                           muxOutVector_11_52_port, A(51) => 
                           muxOutVector_11_51_port, A(50) => 
                           muxOutVector_11_50_port, A(49) => 
                           muxOutVector_11_49_port, A(48) => 
                           muxOutVector_11_48_port, A(47) => 
                           muxOutVector_11_47_port, A(46) => 
                           muxOutVector_11_46_port, A(45) => 
                           muxOutVector_11_45_port, A(44) => 
                           muxOutVector_11_44_port, A(43) => 
                           muxOutVector_11_43_port, A(42) => 
                           muxOutVector_11_42_port, A(41) => 
                           muxOutVector_11_41_port, A(40) => 
                           muxOutVector_11_40_port, A(39) => 
                           muxOutVector_11_39_port, A(38) => 
                           muxOutVector_11_38_port, A(37) => 
                           muxOutVector_11_37_port, A(36) => 
                           muxOutVector_11_36_port, A(35) => 
                           muxOutVector_11_35_port, A(34) => 
                           muxOutVector_11_34_port, A(33) => 
                           muxOutVector_11_33_port, A(32) => 
                           muxOutVector_11_32_port, A(31) => 
                           muxOutVector_11_31_port, A(30) => 
                           muxOutVector_11_30_port, A(29) => 
                           muxOutVector_11_29_port, A(28) => 
                           muxOutVector_11_28_port, A(27) => 
                           muxOutVector_11_27_port, A(26) => 
                           muxOutVector_11_26_port, A(25) => 
                           muxOutVector_11_25_port, A(24) => 
                           muxOutVector_11_24_port, A(23) => 
                           muxOutVector_11_23_port, A(22) => 
                           muxOutVector_11_22_port, A(21) => 
                           muxOutVector_11_21_port, A(20) => 
                           muxOutVector_11_20_port, A(19) => 
                           muxOutVector_11_19_port, A(18) => 
                           muxOutVector_11_18_port, A(17) => 
                           muxOutVector_11_17_port, A(16) => 
                           muxOutVector_11_16_port, A(15) => 
                           muxOutVector_11_15_port, A(14) => 
                           muxOutVector_11_14_port, A(13) => 
                           muxOutVector_11_13_port, A(12) => 
                           muxOutVector_11_12_port, A(11) => 
                           muxOutVector_11_11_port, A(10) => 
                           muxOutVector_11_10_port, A(9) => 
                           muxOutVector_11_9_port, A(8) => 
                           muxOutVector_11_8_port, A(7) => 
                           muxOutVector_11_7_port, A(6) => 
                           muxOutVector_11_6_port, A(5) => 
                           muxOutVector_11_5_port, A(4) => 
                           muxOutVector_11_4_port, A(3) => 
                           muxOutVector_11_3_port, A(2) => 
                           muxOutVector_11_2_port, A(1) => 
                           muxOutVector_11_1_port, A(0) => 
                           muxOutVector_11_0_port, B(63) => 
                           sumVector_10_63_port, B(62) => sumVector_10_62_port,
                           B(61) => sumVector_10_61_port, B(60) => 
                           sumVector_10_60_port, B(59) => sumVector_10_59_port,
                           B(58) => sumVector_10_58_port, B(57) => 
                           sumVector_10_57_port, B(56) => sumVector_10_56_port,
                           B(55) => sumVector_10_55_port, B(54) => 
                           sumVector_10_54_port, B(53) => sumVector_10_53_port,
                           B(52) => sumVector_10_52_port, B(51) => 
                           sumVector_10_51_port, B(50) => sumVector_10_50_port,
                           B(49) => sumVector_10_49_port, B(48) => 
                           sumVector_10_48_port, B(47) => sumVector_10_47_port,
                           B(46) => sumVector_10_46_port, B(45) => 
                           sumVector_10_45_port, B(44) => sumVector_10_44_port,
                           B(43) => sumVector_10_43_port, B(42) => 
                           sumVector_10_42_port, B(41) => sumVector_10_41_port,
                           B(40) => sumVector_10_40_port, B(39) => 
                           sumVector_10_39_port, B(38) => sumVector_10_38_port,
                           B(37) => sumVector_10_37_port, B(36) => 
                           sumVector_10_36_port, B(35) => sumVector_10_35_port,
                           B(34) => sumVector_10_34_port, B(33) => 
                           sumVector_10_33_port, B(32) => sumVector_10_32_port,
                           B(31) => sumVector_10_31_port, B(30) => 
                           sumVector_10_30_port, B(29) => sumVector_10_29_port,
                           B(28) => sumVector_10_28_port, B(27) => 
                           sumVector_10_27_port, B(26) => sumVector_10_26_port,
                           B(25) => sumVector_10_25_port, B(24) => 
                           sumVector_10_24_port, B(23) => sumVector_10_23_port,
                           B(22) => sumVector_10_22_port, B(21) => 
                           sumVector_10_21_port, B(20) => sumVector_10_20_port,
                           B(19) => sumVector_10_19_port, B(18) => 
                           sumVector_10_18_port, B(17) => sumVector_10_17_port,
                           B(16) => sumVector_10_16_port, B(15) => 
                           sumVector_10_15_port, B(14) => sumVector_10_14_port,
                           B(13) => sumVector_10_13_port, B(12) => 
                           sumVector_10_12_port, B(11) => sumVector_10_11_port,
                           B(10) => sumVector_10_10_port, B(9) => 
                           sumVector_10_9_port, B(8) => sumVector_10_8_port, 
                           B(7) => sumVector_10_7_port, B(6) => 
                           sumVector_10_6_port, B(5) => sumVector_10_5_port, 
                           B(4) => sumVector_10_4_port, B(3) => 
                           sumVector_10_3_port, B(2) => sumVector_10_2_port, 
                           B(1) => sumVector_10_1_port, B(0) => 
                           sumVector_10_0_port, Ci => X_Logic0_port, S(63) => 
                           sumVector_11_63_port, S(62) => sumVector_11_62_port,
                           S(61) => sumVector_11_61_port, S(60) => 
                           sumVector_11_60_port, S(59) => sumVector_11_59_port,
                           S(58) => sumVector_11_58_port, S(57) => 
                           sumVector_11_57_port, S(56) => sumVector_11_56_port,
                           S(55) => sumVector_11_55_port, S(54) => 
                           sumVector_11_54_port, S(53) => sumVector_11_53_port,
                           S(52) => sumVector_11_52_port, S(51) => 
                           sumVector_11_51_port, S(50) => sumVector_11_50_port,
                           S(49) => sumVector_11_49_port, S(48) => 
                           sumVector_11_48_port, S(47) => sumVector_11_47_port,
                           S(46) => sumVector_11_46_port, S(45) => 
                           sumVector_11_45_port, S(44) => sumVector_11_44_port,
                           S(43) => sumVector_11_43_port, S(42) => 
                           sumVector_11_42_port, S(41) => sumVector_11_41_port,
                           S(40) => sumVector_11_40_port, S(39) => 
                           sumVector_11_39_port, S(38) => sumVector_11_38_port,
                           S(37) => sumVector_11_37_port, S(36) => 
                           sumVector_11_36_port, S(35) => sumVector_11_35_port,
                           S(34) => sumVector_11_34_port, S(33) => 
                           sumVector_11_33_port, S(32) => sumVector_11_32_port,
                           S(31) => sumVector_11_31_port, S(30) => 
                           sumVector_11_30_port, S(29) => sumVector_11_29_port,
                           S(28) => sumVector_11_28_port, S(27) => 
                           sumVector_11_27_port, S(26) => sumVector_11_26_port,
                           S(25) => sumVector_11_25_port, S(24) => 
                           sumVector_11_24_port, S(23) => sumVector_11_23_port,
                           S(22) => sumVector_11_22_port, S(21) => 
                           sumVector_11_21_port, S(20) => sumVector_11_20_port,
                           S(19) => sumVector_11_19_port, S(18) => 
                           sumVector_11_18_port, S(17) => sumVector_11_17_port,
                           S(16) => sumVector_11_16_port, S(15) => 
                           sumVector_11_15_port, S(14) => sumVector_11_14_port,
                           S(13) => sumVector_11_13_port, S(12) => 
                           sumVector_11_12_port, S(11) => sumVector_11_11_port,
                           S(10) => sumVector_11_10_port, S(9) => 
                           sumVector_11_9_port, S(8) => sumVector_11_8_port, 
                           S(7) => sumVector_11_7_port, S(6) => 
                           sumVector_11_6_port, S(5) => sumVector_11_5_port, 
                           S(4) => sumVector_11_4_port, S(3) => 
                           sumVector_11_3_port, S(2) => sumVector_11_2_port, 
                           S(1) => sumVector_11_1_port, S(0) => 
                           sumVector_11_0_port, Co => n_1046);
   mux_11 : MUX_5TO1_NBIT64_5 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n122, A1(62) => n122, 
                           A1(61) => n121, A1(60) => n121, A1(59) => n121, 
                           A1(58) => n121, A1(57) => n121, A1(56) => n121, 
                           A1(55) => n121, A1(54) => n121, A1(53) => n121, 
                           A1(52) => n374, A1(51) => n367, A1(50) => n360, 
                           A1(49) => n353, A1(48) => n346, A1(47) => n339, 
                           A1(46) => n332, A1(45) => n325, A1(44) => n318, 
                           A1(43) => n311, A1(42) => n304, A1(41) => n297, 
                           A1(40) => n290, A1(39) => n283, A1(38) => n276, 
                           A1(37) => n269, A1(36) => n262, A1(35) => n255, 
                           A1(34) => n248, A1(33) => n241, A1(32) => n234, 
                           A1(31) => n227, A1(30) => n220, A1(29) => n213, 
                           A1(28) => n206, A1(27) => n199, A1(26) => n192, 
                           A1(25) => n186, A1(24) => n182, A1(23) => n176, 
                           A1(22) => A(0), A1(21) => X_Logic0_port, A1(20) => 
                           X_Logic0_port, A1(19) => X_Logic0_port, A1(18) => 
                           X_Logic0_port, A1(17) => X_Logic0_port, A1(16) => 
                           X_Logic0_port, A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(63) => n521, A2(62) => n521, 
                           A2(61) => n520, A2(60) => n520, A2(59) => n520, 
                           A2(58) => n520, A2(57) => n520, A2(56) => n520, 
                           A2(55) => n520, A2(54) => n520, A2(53) => n493, 
                           A2(52) => n489, A2(51) => n485, A2(50) => n481, 
                           A2(49) => n477, A2(48) => n473, A2(47) => n469, 
                           A2(46) => n465, A2(45) => n461, A2(44) => n457, 
                           A2(43) => n453, A2(42) => n449, A2(41) => n445, 
                           A2(40) => n441, A2(39) => n437, A2(38) => n433, 
                           A2(37) => n430, A2(36) => n426, A2(35) => n423, 
                           A2(34) => n420, A2(33) => n416, A2(32) => n412, 
                           A2(31) => n409, A2(30) => n405, A2(29) => n401, 
                           A2(28) => n105, A2(27) => n394, A2(26) => n392, 
                           A2(25) => n389, A2(24) => n387, A2(23) => n383, 
                           A2(22) => n168, A2(21) => X_Logic0_port, A2(20) => 
                           X_Logic0_port, A2(19) => X_Logic0_port, A2(18) => 
                           X_Logic0_port, A2(17) => X_Logic0_port, A2(16) => 
                           X_Logic0_port, A2(15) => X_Logic0_port, A2(14) => 
                           X_Logic0_port, A2(13) => X_Logic0_port, A2(12) => 
                           X_Logic0_port, A2(11) => X_Logic0_port, A2(10) => 
                           X_Logic0_port, A2(9) => X_Logic0_port, A2(8) => 
                           X_Logic0_port, A2(7) => X_Logic0_port, A2(6) => 
                           X_Logic0_port, A2(5) => X_Logic0_port, A2(4) => 
                           X_Logic0_port, A2(3) => X_Logic0_port, A2(2) => 
                           X_Logic0_port, A2(1) => X_Logic0_port, A2(0) => 
                           X_Logic0_port, A3(63) => n153, A3(62) => n153, 
                           A3(61) => n153, A3(60) => n153, A3(59) => n153, 
                           A3(58) => n153, A3(57) => n153, A3(56) => n153, 
                           A3(55) => n153, A3(54) => n153, A3(53) => n377, 
                           A3(52) => n370, A3(51) => n363, A3(50) => n356, 
                           A3(49) => n349, A3(48) => n342, A3(47) => n335, 
                           A3(46) => n328, A3(45) => n321, A3(44) => n314, 
                           A3(43) => n307, A3(42) => n300, A3(41) => n293, 
                           A3(40) => n286, A3(39) => n279, A3(38) => n272, 
                           A3(37) => n265, A3(36) => n258, A3(35) => n251, 
                           A3(34) => n244, A3(33) => n237, A3(32) => n230, 
                           A3(31) => n223, A3(30) => n216, A3(29) => n209, 
                           A3(28) => n202, A3(27) => n195, A3(26) => n186, 
                           A3(25) => n182, A3(24) => n103, A3(23) => A(0), 
                           A3(22) => X_Logic0_port, A3(21) => X_Logic0_port, 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n506, A4(62) => 
                           n506, A4(61) => n506, A4(60) => n506, A4(59) => n505
                           , A4(58) => n505, A4(57) => n505, A4(56) => n505, 
                           A4(55) => n505, A4(54) => n493, A4(53) => n489, 
                           A4(52) => n485, A4(51) => n481, A4(50) => n477, 
                           A4(49) => n473, A4(48) => n469, A4(47) => n465, 
                           A4(46) => n461, A4(45) => n457, A4(44) => n453, 
                           A4(43) => n449, A4(42) => n445, A4(41) => n441, 
                           A4(40) => n437, A4(39) => n433, A4(38) => n430, 
                           A4(37) => n426, A4(36) => n423, A4(35) => n420, 
                           A4(34) => n416, A4(33) => n412, A4(32) => n409, 
                           A4(31) => n405, A4(30) => n401, A4(29) => n104, 
                           A4(28) => n394, A4(27) => n392, A4(26) => n100, 
                           A4(25) => n387, A4(24) => n99, A4(23) => n168, 
                           A4(22) => X_Logic0_port, A4(21) => X_Logic0_port, 
                           A4(20) => X_Logic0_port, A4(19) => X_Logic0_port, 
                           A4(18) => X_Logic0_port, A4(17) => X_Logic0_port, 
                           A4(16) => X_Logic0_port, A4(15) => X_Logic0_port, 
                           A4(14) => X_Logic0_port, A4(13) => X_Logic0_port, 
                           A4(12) => X_Logic0_port, A4(11) => X_Logic0_port, 
                           A4(10) => X_Logic0_port, A4(9) => X_Logic0_port, 
                           A4(8) => X_Logic0_port, A4(7) => X_Logic0_port, 
                           A4(6) => X_Logic0_port, A4(5) => X_Logic0_port, 
                           A4(4) => X_Logic0_port, A4(3) => X_Logic0_port, 
                           A4(2) => X_Logic0_port, A4(1) => X_Logic0_port, 
                           A4(0) => X_Logic0_port, sel(2) => 
                           selVector_11_2_port, sel(1) => selVector_11_1_port, 
                           sel(0) => selVector_11_0_port, O(63) => 
                           muxOutVector_11_63_port, O(62) => 
                           muxOutVector_11_62_port, O(61) => 
                           muxOutVector_11_61_port, O(60) => 
                           muxOutVector_11_60_port, O(59) => 
                           muxOutVector_11_59_port, O(58) => 
                           muxOutVector_11_58_port, O(57) => 
                           muxOutVector_11_57_port, O(56) => 
                           muxOutVector_11_56_port, O(55) => 
                           muxOutVector_11_55_port, O(54) => 
                           muxOutVector_11_54_port, O(53) => 
                           muxOutVector_11_53_port, O(52) => 
                           muxOutVector_11_52_port, O(51) => 
                           muxOutVector_11_51_port, O(50) => 
                           muxOutVector_11_50_port, O(49) => 
                           muxOutVector_11_49_port, O(48) => 
                           muxOutVector_11_48_port, O(47) => 
                           muxOutVector_11_47_port, O(46) => 
                           muxOutVector_11_46_port, O(45) => 
                           muxOutVector_11_45_port, O(44) => 
                           muxOutVector_11_44_port, O(43) => 
                           muxOutVector_11_43_port, O(42) => 
                           muxOutVector_11_42_port, O(41) => 
                           muxOutVector_11_41_port, O(40) => 
                           muxOutVector_11_40_port, O(39) => 
                           muxOutVector_11_39_port, O(38) => 
                           muxOutVector_11_38_port, O(37) => 
                           muxOutVector_11_37_port, O(36) => 
                           muxOutVector_11_36_port, O(35) => 
                           muxOutVector_11_35_port, O(34) => 
                           muxOutVector_11_34_port, O(33) => 
                           muxOutVector_11_33_port, O(32) => 
                           muxOutVector_11_32_port, O(31) => 
                           muxOutVector_11_31_port, O(30) => 
                           muxOutVector_11_30_port, O(29) => 
                           muxOutVector_11_29_port, O(28) => 
                           muxOutVector_11_28_port, O(27) => 
                           muxOutVector_11_27_port, O(26) => 
                           muxOutVector_11_26_port, O(25) => 
                           muxOutVector_11_25_port, O(24) => 
                           muxOutVector_11_24_port, O(23) => 
                           muxOutVector_11_23_port, O(22) => 
                           muxOutVector_11_22_port, O(21) => 
                           muxOutVector_11_21_port, O(20) => 
                           muxOutVector_11_20_port, O(19) => 
                           muxOutVector_11_19_port, O(18) => 
                           muxOutVector_11_18_port, O(17) => 
                           muxOutVector_11_17_port, O(16) => 
                           muxOutVector_11_16_port, O(15) => 
                           muxOutVector_11_15_port, O(14) => 
                           muxOutVector_11_14_port, O(13) => 
                           muxOutVector_11_13_port, O(12) => 
                           muxOutVector_11_12_port, O(11) => 
                           muxOutVector_11_11_port, O(10) => 
                           muxOutVector_11_10_port, O(9) => 
                           muxOutVector_11_9_port, O(8) => 
                           muxOutVector_11_8_port, O(7) => 
                           muxOutVector_11_7_port, O(6) => 
                           muxOutVector_11_6_port, O(5) => 
                           muxOutVector_11_5_port, O(4) => 
                           muxOutVector_11_4_port, O(3) => 
                           muxOutVector_11_3_port, O(2) => 
                           muxOutVector_11_2_port, O(1) => 
                           muxOutVector_11_1_port, O(0) => 
                           muxOutVector_11_0_port);
   eb_12 : BE_BLOCK_4 port map( b(2) => B(25), b(1) => B(24), b(0) => B(23), 
                           sel(2) => selVector_12_2_port, sel(1) => 
                           selVector_12_1_port, sel(0) => selVector_12_0_port);
   sum_12 : RCA_NBIT64_4 port map( A(63) => muxOutVector_12_63_port, A(62) => 
                           muxOutVector_12_62_port, A(61) => 
                           muxOutVector_12_61_port, A(60) => 
                           muxOutVector_12_60_port, A(59) => 
                           muxOutVector_12_59_port, A(58) => 
                           muxOutVector_12_58_port, A(57) => 
                           muxOutVector_12_57_port, A(56) => 
                           muxOutVector_12_56_port, A(55) => 
                           muxOutVector_12_55_port, A(54) => 
                           muxOutVector_12_54_port, A(53) => 
                           muxOutVector_12_53_port, A(52) => 
                           muxOutVector_12_52_port, A(51) => 
                           muxOutVector_12_51_port, A(50) => 
                           muxOutVector_12_50_port, A(49) => 
                           muxOutVector_12_49_port, A(48) => 
                           muxOutVector_12_48_port, A(47) => 
                           muxOutVector_12_47_port, A(46) => 
                           muxOutVector_12_46_port, A(45) => 
                           muxOutVector_12_45_port, A(44) => 
                           muxOutVector_12_44_port, A(43) => 
                           muxOutVector_12_43_port, A(42) => 
                           muxOutVector_12_42_port, A(41) => 
                           muxOutVector_12_41_port, A(40) => 
                           muxOutVector_12_40_port, A(39) => 
                           muxOutVector_12_39_port, A(38) => 
                           muxOutVector_12_38_port, A(37) => 
                           muxOutVector_12_37_port, A(36) => 
                           muxOutVector_12_36_port, A(35) => 
                           muxOutVector_12_35_port, A(34) => 
                           muxOutVector_12_34_port, A(33) => 
                           muxOutVector_12_33_port, A(32) => 
                           muxOutVector_12_32_port, A(31) => 
                           muxOutVector_12_31_port, A(30) => 
                           muxOutVector_12_30_port, A(29) => 
                           muxOutVector_12_29_port, A(28) => 
                           muxOutVector_12_28_port, A(27) => 
                           muxOutVector_12_27_port, A(26) => 
                           muxOutVector_12_26_port, A(25) => 
                           muxOutVector_12_25_port, A(24) => 
                           muxOutVector_12_24_port, A(23) => 
                           muxOutVector_12_23_port, A(22) => 
                           muxOutVector_12_22_port, A(21) => 
                           muxOutVector_12_21_port, A(20) => 
                           muxOutVector_12_20_port, A(19) => 
                           muxOutVector_12_19_port, A(18) => 
                           muxOutVector_12_18_port, A(17) => 
                           muxOutVector_12_17_port, A(16) => 
                           muxOutVector_12_16_port, A(15) => 
                           muxOutVector_12_15_port, A(14) => 
                           muxOutVector_12_14_port, A(13) => 
                           muxOutVector_12_13_port, A(12) => 
                           muxOutVector_12_12_port, A(11) => 
                           muxOutVector_12_11_port, A(10) => 
                           muxOutVector_12_10_port, A(9) => 
                           muxOutVector_12_9_port, A(8) => 
                           muxOutVector_12_8_port, A(7) => 
                           muxOutVector_12_7_port, A(6) => 
                           muxOutVector_12_6_port, A(5) => 
                           muxOutVector_12_5_port, A(4) => 
                           muxOutVector_12_4_port, A(3) => 
                           muxOutVector_12_3_port, A(2) => 
                           muxOutVector_12_2_port, A(1) => 
                           muxOutVector_12_1_port, A(0) => 
                           muxOutVector_12_0_port, B(63) => 
                           sumVector_11_63_port, B(62) => sumVector_11_62_port,
                           B(61) => sumVector_11_61_port, B(60) => 
                           sumVector_11_60_port, B(59) => sumVector_11_59_port,
                           B(58) => sumVector_11_58_port, B(57) => 
                           sumVector_11_57_port, B(56) => sumVector_11_56_port,
                           B(55) => sumVector_11_55_port, B(54) => 
                           sumVector_11_54_port, B(53) => sumVector_11_53_port,
                           B(52) => sumVector_11_52_port, B(51) => 
                           sumVector_11_51_port, B(50) => sumVector_11_50_port,
                           B(49) => sumVector_11_49_port, B(48) => 
                           sumVector_11_48_port, B(47) => sumVector_11_47_port,
                           B(46) => sumVector_11_46_port, B(45) => 
                           sumVector_11_45_port, B(44) => sumVector_11_44_port,
                           B(43) => sumVector_11_43_port, B(42) => 
                           sumVector_11_42_port, B(41) => sumVector_11_41_port,
                           B(40) => sumVector_11_40_port, B(39) => 
                           sumVector_11_39_port, B(38) => sumVector_11_38_port,
                           B(37) => sumVector_11_37_port, B(36) => 
                           sumVector_11_36_port, B(35) => sumVector_11_35_port,
                           B(34) => sumVector_11_34_port, B(33) => 
                           sumVector_11_33_port, B(32) => sumVector_11_32_port,
                           B(31) => sumVector_11_31_port, B(30) => 
                           sumVector_11_30_port, B(29) => sumVector_11_29_port,
                           B(28) => sumVector_11_28_port, B(27) => 
                           sumVector_11_27_port, B(26) => sumVector_11_26_port,
                           B(25) => sumVector_11_25_port, B(24) => 
                           sumVector_11_24_port, B(23) => sumVector_11_23_port,
                           B(22) => sumVector_11_22_port, B(21) => 
                           sumVector_11_21_port, B(20) => sumVector_11_20_port,
                           B(19) => sumVector_11_19_port, B(18) => 
                           sumVector_11_18_port, B(17) => sumVector_11_17_port,
                           B(16) => sumVector_11_16_port, B(15) => 
                           sumVector_11_15_port, B(14) => sumVector_11_14_port,
                           B(13) => sumVector_11_13_port, B(12) => 
                           sumVector_11_12_port, B(11) => sumVector_11_11_port,
                           B(10) => sumVector_11_10_port, B(9) => 
                           sumVector_11_9_port, B(8) => sumVector_11_8_port, 
                           B(7) => sumVector_11_7_port, B(6) => 
                           sumVector_11_6_port, B(5) => sumVector_11_5_port, 
                           B(4) => sumVector_11_4_port, B(3) => 
                           sumVector_11_3_port, B(2) => sumVector_11_2_port, 
                           B(1) => sumVector_11_1_port, B(0) => 
                           sumVector_11_0_port, Ci => X_Logic0_port, S(63) => 
                           sumVector_12_63_port, S(62) => sumVector_12_62_port,
                           S(61) => sumVector_12_61_port, S(60) => 
                           sumVector_12_60_port, S(59) => sumVector_12_59_port,
                           S(58) => sumVector_12_58_port, S(57) => 
                           sumVector_12_57_port, S(56) => sumVector_12_56_port,
                           S(55) => sumVector_12_55_port, S(54) => 
                           sumVector_12_54_port, S(53) => sumVector_12_53_port,
                           S(52) => sumVector_12_52_port, S(51) => 
                           sumVector_12_51_port, S(50) => sumVector_12_50_port,
                           S(49) => sumVector_12_49_port, S(48) => 
                           sumVector_12_48_port, S(47) => sumVector_12_47_port,
                           S(46) => sumVector_12_46_port, S(45) => 
                           sumVector_12_45_port, S(44) => sumVector_12_44_port,
                           S(43) => sumVector_12_43_port, S(42) => 
                           sumVector_12_42_port, S(41) => sumVector_12_41_port,
                           S(40) => sumVector_12_40_port, S(39) => 
                           sumVector_12_39_port, S(38) => sumVector_12_38_port,
                           S(37) => sumVector_12_37_port, S(36) => 
                           sumVector_12_36_port, S(35) => sumVector_12_35_port,
                           S(34) => sumVector_12_34_port, S(33) => 
                           sumVector_12_33_port, S(32) => sumVector_12_32_port,
                           S(31) => sumVector_12_31_port, S(30) => 
                           sumVector_12_30_port, S(29) => sumVector_12_29_port,
                           S(28) => sumVector_12_28_port, S(27) => 
                           sumVector_12_27_port, S(26) => sumVector_12_26_port,
                           S(25) => sumVector_12_25_port, S(24) => 
                           sumVector_12_24_port, S(23) => sumVector_12_23_port,
                           S(22) => sumVector_12_22_port, S(21) => 
                           sumVector_12_21_port, S(20) => sumVector_12_20_port,
                           S(19) => sumVector_12_19_port, S(18) => 
                           sumVector_12_18_port, S(17) => sumVector_12_17_port,
                           S(16) => sumVector_12_16_port, S(15) => 
                           sumVector_12_15_port, S(14) => sumVector_12_14_port,
                           S(13) => sumVector_12_13_port, S(12) => 
                           sumVector_12_12_port, S(11) => sumVector_12_11_port,
                           S(10) => sumVector_12_10_port, S(9) => 
                           sumVector_12_9_port, S(8) => sumVector_12_8_port, 
                           S(7) => sumVector_12_7_port, S(6) => 
                           sumVector_12_6_port, S(5) => sumVector_12_5_port, 
                           S(4) => sumVector_12_4_port, S(3) => 
                           sumVector_12_3_port, S(2) => sumVector_12_2_port, 
                           S(1) => sumVector_12_1_port, S(0) => 
                           sumVector_12_0_port, Co => n_1047);
   mux_12 : MUX_5TO1_NBIT64_4 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n122, A1(62) => n122, 
                           A1(61) => n122, A1(60) => n125, A1(59) => n122, 
                           A1(58) => n122, A1(57) => n122, A1(56) => n122, 
                           A1(55) => n122, A1(54) => n376, A1(53) => n369, 
                           A1(52) => n362, A1(51) => n355, A1(50) => n348, 
                           A1(49) => n341, A1(48) => n334, A1(47) => n327, 
                           A1(46) => n320, A1(45) => n313, A1(44) => n306, 
                           A1(43) => n299, A1(42) => n292, A1(41) => n285, 
                           A1(40) => n278, A1(39) => n271, A1(38) => n264, 
                           A1(37) => n257, A1(36) => n250, A1(35) => n243, 
                           A1(34) => n236, A1(33) => n229, A1(32) => n222, 
                           A1(31) => n215, A1(30) => n208, A1(29) => n201, 
                           A1(28) => n194, A1(27) => n186, A1(26) => n182, 
                           A1(25) => n176, A1(24) => A(0), A1(23) => 
                           X_Logic0_port, A1(22) => X_Logic0_port, A1(21) => 
                           X_Logic0_port, A1(20) => X_Logic0_port, A1(19) => 
                           X_Logic0_port, A1(18) => X_Logic0_port, A1(17) => 
                           X_Logic0_port, A1(16) => X_Logic0_port, A1(15) => 
                           X_Logic0_port, A1(14) => X_Logic0_port, A1(13) => 
                           X_Logic0_port, A1(12) => X_Logic0_port, A1(11) => 
                           X_Logic0_port, A1(10) => X_Logic0_port, A1(9) => 
                           X_Logic0_port, A1(8) => X_Logic0_port, A1(7) => 
                           X_Logic0_port, A1(6) => X_Logic0_port, A1(5) => 
                           X_Logic0_port, A1(4) => X_Logic0_port, A1(3) => 
                           X_Logic0_port, A1(2) => X_Logic0_port, A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n522, A2(62) => n522, A2(61) => n522, A2(60) => n522
                           , A2(59) => n522, A2(58) => n522, A2(57) => n521, 
                           A2(56) => n521, A2(55) => n493, A2(54) => n489, 
                           A2(53) => n485, A2(52) => n481, A2(51) => n477, 
                           A2(50) => n473, A2(49) => n469, A2(48) => n465, 
                           A2(47) => n461, A2(46) => n457, A2(45) => n453, 
                           A2(44) => n449, A2(43) => n445, A2(42) => n441, 
                           A2(41) => n437, A2(40) => n433, A2(39) => n430, 
                           A2(38) => n426, A2(37) => n423, A2(36) => n420, 
                           A2(35) => n416, A2(34) => n412, A2(33) => n409, 
                           A2(32) => n405, A2(31) => n401, A2(30) => n398, 
                           A2(29) => n396, A2(28) => n392, A2(27) => n101, 
                           A2(26) => n387, A2(25) => n99, A2(24) => n168, 
                           A2(23) => X_Logic0_port, A2(22) => X_Logic0_port, 
                           A2(21) => X_Logic0_port, A2(20) => X_Logic0_port, 
                           A2(19) => X_Logic0_port, A2(18) => X_Logic0_port, 
                           A2(17) => X_Logic0_port, A2(16) => X_Logic0_port, 
                           A2(15) => X_Logic0_port, A2(14) => X_Logic0_port, 
                           A2(13) => X_Logic0_port, A2(12) => X_Logic0_port, 
                           A2(11) => X_Logic0_port, A2(10) => X_Logic0_port, 
                           A2(9) => X_Logic0_port, A2(8) => X_Logic0_port, 
                           A2(7) => X_Logic0_port, A2(6) => X_Logic0_port, 
                           A2(5) => X_Logic0_port, A2(4) => X_Logic0_port, 
                           A2(3) => X_Logic0_port, A2(2) => X_Logic0_port, 
                           A2(1) => X_Logic0_port, A2(0) => X_Logic0_port, 
                           A3(63) => n152, A3(62) => n152, A3(61) => n152, 
                           A3(60) => n152, A3(59) => n152, A3(58) => n152, 
                           A3(57) => n152, A3(56) => n152, A3(55) => n378, 
                           A3(54) => n371, A3(53) => n364, A3(52) => n357, 
                           A3(51) => n350, A3(50) => n343, A3(49) => n336, 
                           A3(48) => n329, A3(47) => n322, A3(46) => n315, 
                           A3(45) => n308, A3(44) => n301, A3(43) => n294, 
                           A3(42) => n287, A3(41) => n280, A3(40) => n273, 
                           A3(39) => n266, A3(38) => n259, A3(37) => n252, 
                           A3(36) => n245, A3(35) => n238, A3(34) => n231, 
                           A3(33) => n224, A3(32) => n217, A3(31) => n210, 
                           A3(30) => n203, A3(29) => n196, A3(28) => n186, 
                           A3(27) => n182, A3(26) => n103, A3(25) => A(0), 
                           A3(24) => X_Logic0_port, A3(23) => X_Logic0_port, 
                           A3(22) => X_Logic0_port, A3(21) => X_Logic0_port, 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n506, A4(62) => 
                           n506, A4(61) => n506, A4(60) => n506, A4(59) => n506
                           , A4(58) => n506, A4(57) => n506, A4(56) => n493, 
                           A4(55) => n489, A4(54) => n485, A4(53) => n481, 
                           A4(52) => n477, A4(51) => n473, A4(50) => n469, 
                           A4(49) => n465, A4(48) => n461, A4(47) => n457, 
                           A4(46) => n453, A4(45) => n449, A4(44) => n445, 
                           A4(43) => n441, A4(42) => n437, A4(41) => n433, 
                           A4(40) => n430, A4(39) => n426, A4(38) => n423, 
                           A4(37) => n420, A4(36) => n416, A4(35) => n412, 
                           A4(34) => n409, A4(33) => n405, A4(32) => n401, 
                           A4(31) => n397, A4(30) => n396, A4(29) => n392, 
                           A4(28) => n388, A4(27) => n387, A4(26) => n99, 
                           A4(25) => n167, A4(24) => X_Logic0_port, A4(23) => 
                           X_Logic0_port, A4(22) => X_Logic0_port, A4(21) => 
                           X_Logic0_port, A4(20) => X_Logic0_port, A4(19) => 
                           X_Logic0_port, A4(18) => X_Logic0_port, A4(17) => 
                           X_Logic0_port, A4(16) => X_Logic0_port, A4(15) => 
                           X_Logic0_port, A4(14) => X_Logic0_port, A4(13) => 
                           X_Logic0_port, A4(12) => X_Logic0_port, A4(11) => 
                           X_Logic0_port, A4(10) => X_Logic0_port, A4(9) => 
                           X_Logic0_port, A4(8) => X_Logic0_port, A4(7) => 
                           X_Logic0_port, A4(6) => X_Logic0_port, A4(5) => 
                           X_Logic0_port, A4(4) => X_Logic0_port, A4(3) => 
                           X_Logic0_port, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_12_2_port, sel(1) => selVector_12_1_port, 
                           sel(0) => selVector_12_0_port, O(63) => 
                           muxOutVector_12_63_port, O(62) => 
                           muxOutVector_12_62_port, O(61) => 
                           muxOutVector_12_61_port, O(60) => 
                           muxOutVector_12_60_port, O(59) => 
                           muxOutVector_12_59_port, O(58) => 
                           muxOutVector_12_58_port, O(57) => 
                           muxOutVector_12_57_port, O(56) => 
                           muxOutVector_12_56_port, O(55) => 
                           muxOutVector_12_55_port, O(54) => 
                           muxOutVector_12_54_port, O(53) => 
                           muxOutVector_12_53_port, O(52) => 
                           muxOutVector_12_52_port, O(51) => 
                           muxOutVector_12_51_port, O(50) => 
                           muxOutVector_12_50_port, O(49) => 
                           muxOutVector_12_49_port, O(48) => 
                           muxOutVector_12_48_port, O(47) => 
                           muxOutVector_12_47_port, O(46) => 
                           muxOutVector_12_46_port, O(45) => 
                           muxOutVector_12_45_port, O(44) => 
                           muxOutVector_12_44_port, O(43) => 
                           muxOutVector_12_43_port, O(42) => 
                           muxOutVector_12_42_port, O(41) => 
                           muxOutVector_12_41_port, O(40) => 
                           muxOutVector_12_40_port, O(39) => 
                           muxOutVector_12_39_port, O(38) => 
                           muxOutVector_12_38_port, O(37) => 
                           muxOutVector_12_37_port, O(36) => 
                           muxOutVector_12_36_port, O(35) => 
                           muxOutVector_12_35_port, O(34) => 
                           muxOutVector_12_34_port, O(33) => 
                           muxOutVector_12_33_port, O(32) => 
                           muxOutVector_12_32_port, O(31) => 
                           muxOutVector_12_31_port, O(30) => 
                           muxOutVector_12_30_port, O(29) => 
                           muxOutVector_12_29_port, O(28) => 
                           muxOutVector_12_28_port, O(27) => 
                           muxOutVector_12_27_port, O(26) => 
                           muxOutVector_12_26_port, O(25) => 
                           muxOutVector_12_25_port, O(24) => 
                           muxOutVector_12_24_port, O(23) => 
                           muxOutVector_12_23_port, O(22) => 
                           muxOutVector_12_22_port, O(21) => 
                           muxOutVector_12_21_port, O(20) => 
                           muxOutVector_12_20_port, O(19) => 
                           muxOutVector_12_19_port, O(18) => 
                           muxOutVector_12_18_port, O(17) => 
                           muxOutVector_12_17_port, O(16) => 
                           muxOutVector_12_16_port, O(15) => 
                           muxOutVector_12_15_port, O(14) => 
                           muxOutVector_12_14_port, O(13) => 
                           muxOutVector_12_13_port, O(12) => 
                           muxOutVector_12_12_port, O(11) => 
                           muxOutVector_12_11_port, O(10) => 
                           muxOutVector_12_10_port, O(9) => 
                           muxOutVector_12_9_port, O(8) => 
                           muxOutVector_12_8_port, O(7) => 
                           muxOutVector_12_7_port, O(6) => 
                           muxOutVector_12_6_port, O(5) => 
                           muxOutVector_12_5_port, O(4) => 
                           muxOutVector_12_4_port, O(3) => 
                           muxOutVector_12_3_port, O(2) => 
                           muxOutVector_12_2_port, O(1) => 
                           muxOutVector_12_1_port, O(0) => 
                           muxOutVector_12_0_port);
   eb_13 : BE_BLOCK_3 port map( b(2) => B(27), b(1) => B(26), b(0) => B(25), 
                           sel(2) => selVector_13_2_port, sel(1) => 
                           selVector_13_1_port, sel(0) => selVector_13_0_port);
   sum_13 : RCA_NBIT64_3 port map( A(63) => muxOutVector_13_63_port, A(62) => 
                           muxOutVector_13_62_port, A(61) => 
                           muxOutVector_13_61_port, A(60) => 
                           muxOutVector_13_60_port, A(59) => 
                           muxOutVector_13_59_port, A(58) => 
                           muxOutVector_13_58_port, A(57) => 
                           muxOutVector_13_57_port, A(56) => 
                           muxOutVector_13_56_port, A(55) => 
                           muxOutVector_13_55_port, A(54) => 
                           muxOutVector_13_54_port, A(53) => 
                           muxOutVector_13_53_port, A(52) => 
                           muxOutVector_13_52_port, A(51) => 
                           muxOutVector_13_51_port, A(50) => 
                           muxOutVector_13_50_port, A(49) => 
                           muxOutVector_13_49_port, A(48) => 
                           muxOutVector_13_48_port, A(47) => 
                           muxOutVector_13_47_port, A(46) => 
                           muxOutVector_13_46_port, A(45) => 
                           muxOutVector_13_45_port, A(44) => 
                           muxOutVector_13_44_port, A(43) => 
                           muxOutVector_13_43_port, A(42) => 
                           muxOutVector_13_42_port, A(41) => 
                           muxOutVector_13_41_port, A(40) => 
                           muxOutVector_13_40_port, A(39) => 
                           muxOutVector_13_39_port, A(38) => 
                           muxOutVector_13_38_port, A(37) => 
                           muxOutVector_13_37_port, A(36) => 
                           muxOutVector_13_36_port, A(35) => 
                           muxOutVector_13_35_port, A(34) => 
                           muxOutVector_13_34_port, A(33) => 
                           muxOutVector_13_33_port, A(32) => 
                           muxOutVector_13_32_port, A(31) => 
                           muxOutVector_13_31_port, A(30) => 
                           muxOutVector_13_30_port, A(29) => 
                           muxOutVector_13_29_port, A(28) => 
                           muxOutVector_13_28_port, A(27) => 
                           muxOutVector_13_27_port, A(26) => 
                           muxOutVector_13_26_port, A(25) => 
                           muxOutVector_13_25_port, A(24) => 
                           muxOutVector_13_24_port, A(23) => 
                           muxOutVector_13_23_port, A(22) => 
                           muxOutVector_13_22_port, A(21) => 
                           muxOutVector_13_21_port, A(20) => 
                           muxOutVector_13_20_port, A(19) => 
                           muxOutVector_13_19_port, A(18) => 
                           muxOutVector_13_18_port, A(17) => 
                           muxOutVector_13_17_port, A(16) => 
                           muxOutVector_13_16_port, A(15) => 
                           muxOutVector_13_15_port, A(14) => 
                           muxOutVector_13_14_port, A(13) => 
                           muxOutVector_13_13_port, A(12) => 
                           muxOutVector_13_12_port, A(11) => 
                           muxOutVector_13_11_port, A(10) => 
                           muxOutVector_13_10_port, A(9) => 
                           muxOutVector_13_9_port, A(8) => 
                           muxOutVector_13_8_port, A(7) => 
                           muxOutVector_13_7_port, A(6) => 
                           muxOutVector_13_6_port, A(5) => 
                           muxOutVector_13_5_port, A(4) => 
                           muxOutVector_13_4_port, A(3) => 
                           muxOutVector_13_3_port, A(2) => 
                           muxOutVector_13_2_port, A(1) => 
                           muxOutVector_13_1_port, A(0) => 
                           muxOutVector_13_0_port, B(63) => 
                           sumVector_12_63_port, B(62) => sumVector_12_62_port,
                           B(61) => sumVector_12_61_port, B(60) => 
                           sumVector_12_60_port, B(59) => sumVector_12_59_port,
                           B(58) => sumVector_12_58_port, B(57) => 
                           sumVector_12_57_port, B(56) => sumVector_12_56_port,
                           B(55) => sumVector_12_55_port, B(54) => 
                           sumVector_12_54_port, B(53) => sumVector_12_53_port,
                           B(52) => sumVector_12_52_port, B(51) => 
                           sumVector_12_51_port, B(50) => sumVector_12_50_port,
                           B(49) => sumVector_12_49_port, B(48) => 
                           sumVector_12_48_port, B(47) => sumVector_12_47_port,
                           B(46) => sumVector_12_46_port, B(45) => 
                           sumVector_12_45_port, B(44) => sumVector_12_44_port,
                           B(43) => sumVector_12_43_port, B(42) => 
                           sumVector_12_42_port, B(41) => sumVector_12_41_port,
                           B(40) => sumVector_12_40_port, B(39) => 
                           sumVector_12_39_port, B(38) => sumVector_12_38_port,
                           B(37) => sumVector_12_37_port, B(36) => 
                           sumVector_12_36_port, B(35) => sumVector_12_35_port,
                           B(34) => sumVector_12_34_port, B(33) => 
                           sumVector_12_33_port, B(32) => sumVector_12_32_port,
                           B(31) => sumVector_12_31_port, B(30) => 
                           sumVector_12_30_port, B(29) => sumVector_12_29_port,
                           B(28) => sumVector_12_28_port, B(27) => 
                           sumVector_12_27_port, B(26) => sumVector_12_26_port,
                           B(25) => sumVector_12_25_port, B(24) => 
                           sumVector_12_24_port, B(23) => sumVector_12_23_port,
                           B(22) => sumVector_12_22_port, B(21) => 
                           sumVector_12_21_port, B(20) => sumVector_12_20_port,
                           B(19) => sumVector_12_19_port, B(18) => 
                           sumVector_12_18_port, B(17) => sumVector_12_17_port,
                           B(16) => sumVector_12_16_port, B(15) => 
                           sumVector_12_15_port, B(14) => sumVector_12_14_port,
                           B(13) => sumVector_12_13_port, B(12) => 
                           sumVector_12_12_port, B(11) => sumVector_12_11_port,
                           B(10) => sumVector_12_10_port, B(9) => 
                           sumVector_12_9_port, B(8) => sumVector_12_8_port, 
                           B(7) => sumVector_12_7_port, B(6) => 
                           sumVector_12_6_port, B(5) => sumVector_12_5_port, 
                           B(4) => sumVector_12_4_port, B(3) => 
                           sumVector_12_3_port, B(2) => sumVector_12_2_port, 
                           B(1) => sumVector_12_1_port, B(0) => 
                           sumVector_12_0_port, Ci => X_Logic0_port, S(63) => 
                           sumVector_13_63_port, S(62) => sumVector_13_62_port,
                           S(61) => sumVector_13_61_port, S(60) => 
                           sumVector_13_60_port, S(59) => sumVector_13_59_port,
                           S(58) => sumVector_13_58_port, S(57) => 
                           sumVector_13_57_port, S(56) => sumVector_13_56_port,
                           S(55) => sumVector_13_55_port, S(54) => 
                           sumVector_13_54_port, S(53) => sumVector_13_53_port,
                           S(52) => sumVector_13_52_port, S(51) => 
                           sumVector_13_51_port, S(50) => sumVector_13_50_port,
                           S(49) => sumVector_13_49_port, S(48) => 
                           sumVector_13_48_port, S(47) => sumVector_13_47_port,
                           S(46) => sumVector_13_46_port, S(45) => 
                           sumVector_13_45_port, S(44) => sumVector_13_44_port,
                           S(43) => sumVector_13_43_port, S(42) => 
                           sumVector_13_42_port, S(41) => sumVector_13_41_port,
                           S(40) => sumVector_13_40_port, S(39) => 
                           sumVector_13_39_port, S(38) => sumVector_13_38_port,
                           S(37) => sumVector_13_37_port, S(36) => 
                           sumVector_13_36_port, S(35) => sumVector_13_35_port,
                           S(34) => sumVector_13_34_port, S(33) => 
                           sumVector_13_33_port, S(32) => sumVector_13_32_port,
                           S(31) => sumVector_13_31_port, S(30) => 
                           sumVector_13_30_port, S(29) => sumVector_13_29_port,
                           S(28) => sumVector_13_28_port, S(27) => 
                           sumVector_13_27_port, S(26) => sumVector_13_26_port,
                           S(25) => sumVector_13_25_port, S(24) => 
                           sumVector_13_24_port, S(23) => sumVector_13_23_port,
                           S(22) => sumVector_13_22_port, S(21) => 
                           sumVector_13_21_port, S(20) => sumVector_13_20_port,
                           S(19) => sumVector_13_19_port, S(18) => 
                           sumVector_13_18_port, S(17) => sumVector_13_17_port,
                           S(16) => sumVector_13_16_port, S(15) => 
                           sumVector_13_15_port, S(14) => sumVector_13_14_port,
                           S(13) => sumVector_13_13_port, S(12) => 
                           sumVector_13_12_port, S(11) => sumVector_13_11_port,
                           S(10) => sumVector_13_10_port, S(9) => 
                           sumVector_13_9_port, S(8) => sumVector_13_8_port, 
                           S(7) => sumVector_13_7_port, S(6) => 
                           sumVector_13_6_port, S(5) => sumVector_13_5_port, 
                           S(4) => sumVector_13_4_port, S(3) => 
                           sumVector_13_3_port, S(2) => sumVector_13_2_port, 
                           S(1) => sumVector_13_1_port, S(0) => 
                           sumVector_13_0_port, Co => n_1048);
   mux_13 : MUX_5TO1_NBIT64_3 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n123, A1(62) => n123, 
                           A1(61) => n123, A1(60) => n123, A1(59) => n123, 
                           A1(58) => n123, A1(57) => n122, A1(56) => n375, 
                           A1(55) => n368, A1(54) => n361, A1(53) => n354, 
                           A1(52) => n347, A1(51) => n340, A1(50) => n333, 
                           A1(49) => n326, A1(48) => n319, A1(47) => n312, 
                           A1(46) => n305, A1(45) => n298, A1(44) => n291, 
                           A1(43) => n284, A1(42) => n277, A1(41) => n270, 
                           A1(40) => n263, A1(39) => n256, A1(38) => n249, 
                           A1(37) => n242, A1(36) => n235, A1(35) => n228, 
                           A1(34) => n221, A1(33) => n214, A1(32) => n207, 
                           A1(31) => n200, A1(30) => n193, A1(29) => n186, 
                           A1(28) => n182, A1(27) => n176, A1(26) => A(0), 
                           A1(25) => X_Logic0_port, A1(24) => X_Logic0_port, 
                           A1(23) => X_Logic0_port, A1(22) => X_Logic0_port, 
                           A1(21) => X_Logic0_port, A1(20) => X_Logic0_port, 
                           A1(19) => X_Logic0_port, A1(18) => X_Logic0_port, 
                           A1(17) => X_Logic0_port, A1(16) => X_Logic0_port, 
                           A1(15) => X_Logic0_port, A1(14) => X_Logic0_port, 
                           A1(13) => X_Logic0_port, A1(12) => X_Logic0_port, 
                           A1(11) => X_Logic0_port, A1(10) => X_Logic0_port, 
                           A1(9) => X_Logic0_port, A1(8) => X_Logic0_port, 
                           A1(7) => X_Logic0_port, A1(6) => X_Logic0_port, 
                           A1(5) => X_Logic0_port, A1(4) => X_Logic0_port, 
                           A1(3) => X_Logic0_port, A1(2) => X_Logic0_port, 
                           A1(1) => X_Logic0_port, A1(0) => X_Logic0_port, 
                           A2(63) => n523, A2(62) => n523, A2(61) => n523, 
                           A2(60) => n523, A2(59) => n523, A2(58) => n522, 
                           A2(57) => n493, A2(56) => n489, A2(55) => n485, 
                           A2(54) => n481, A2(53) => n477, A2(52) => n473, 
                           A2(51) => n469, A2(50) => n465, A2(49) => n461, 
                           A2(48) => n457, A2(47) => n453, A2(46) => n449, 
                           A2(45) => n445, A2(44) => n441, A2(43) => n437, 
                           A2(42) => n433, A2(41) => n430, A2(40) => n426, 
                           A2(39) => n423, A2(38) => n420, A2(37) => n416, 
                           A2(36) => n412, A2(35) => n409, A2(34) => n405, 
                           A2(33) => n401, A2(32) => n105, A2(31) => n394, 
                           A2(30) => n392, A2(29) => n100, A2(28) => n387, 
                           A2(27) => n383, A2(26) => n168, A2(25) => 
                           X_Logic0_port, A2(24) => X_Logic0_port, A2(23) => 
                           X_Logic0_port, A2(22) => X_Logic0_port, A2(21) => 
                           X_Logic0_port, A2(20) => X_Logic0_port, A2(19) => 
                           X_Logic0_port, A2(18) => X_Logic0_port, A2(17) => 
                           X_Logic0_port, A2(16) => X_Logic0_port, A2(15) => 
                           X_Logic0_port, A2(14) => X_Logic0_port, A2(13) => 
                           X_Logic0_port, A2(12) => X_Logic0_port, A2(11) => 
                           X_Logic0_port, A2(10) => X_Logic0_port, A2(9) => 
                           X_Logic0_port, A2(8) => X_Logic0_port, A2(7) => 
                           X_Logic0_port, A2(6) => X_Logic0_port, A2(5) => 
                           X_Logic0_port, A2(4) => X_Logic0_port, A2(3) => 
                           X_Logic0_port, A2(2) => X_Logic0_port, A2(1) => 
                           X_Logic0_port, A2(0) => X_Logic0_port, A3(63) => 
                           n151, A3(62) => n151, A3(61) => n152, A3(60) => n152
                           , A3(59) => n152, A3(58) => n152, A3(57) => n375, 
                           A3(56) => n368, A3(55) => n361, A3(54) => n354, 
                           A3(53) => n347, A3(52) => n340, A3(51) => n333, 
                           A3(50) => n326, A3(49) => n319, A3(48) => n312, 
                           A3(47) => n305, A3(46) => n298, A3(45) => n291, 
                           A3(44) => n284, A3(43) => n277, A3(42) => n270, 
                           A3(41) => n263, A3(40) => n256, A3(39) => n249, 
                           A3(38) => n242, A3(37) => n235, A3(36) => n228, 
                           A3(35) => n221, A3(34) => n214, A3(33) => n207, 
                           A3(32) => n200, A3(31) => n193, A3(30) => n186, 
                           A3(29) => n182, A3(28) => n103, A3(27) => A(0), 
                           A3(26) => X_Logic0_port, A3(25) => X_Logic0_port, 
                           A3(24) => X_Logic0_port, A3(23) => X_Logic0_port, 
                           A3(22) => X_Logic0_port, A3(21) => X_Logic0_port, 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n507, A4(62) => 
                           n507, A4(61) => n507, A4(60) => n507, A4(59) => n506
                           , A4(58) => n492, A4(57) => n488, A4(56) => n484, 
                           A4(55) => n480, A4(54) => n476, A4(53) => n472, 
                           A4(52) => n468, A4(51) => n464, A4(50) => n460, 
                           A4(49) => n456, A4(48) => n452, A4(47) => n448, 
                           A4(46) => n444, A4(45) => n440, A4(44) => n436, 
                           A4(43) => n432, A4(42) => n429, A4(41) => n425, 
                           A4(40) => n422, A4(39) => n419, A4(38) => n415, 
                           A4(37) => n411, A4(36) => n408, A4(35) => n404, 
                           A4(34) => n400, A4(33) => n104, A4(32) => n396, 
                           A4(31) => n391, A4(30) => n389, A4(29) => n386, 
                           A4(28) => n385, A4(27) => n167, A4(26) => 
                           X_Logic0_port, A4(25) => X_Logic0_port, A4(24) => 
                           X_Logic0_port, A4(23) => X_Logic0_port, A4(22) => 
                           X_Logic0_port, A4(21) => X_Logic0_port, A4(20) => 
                           X_Logic0_port, A4(19) => X_Logic0_port, A4(18) => 
                           X_Logic0_port, A4(17) => X_Logic0_port, A4(16) => 
                           X_Logic0_port, A4(15) => X_Logic0_port, A4(14) => 
                           X_Logic0_port, A4(13) => X_Logic0_port, A4(12) => 
                           X_Logic0_port, A4(11) => X_Logic0_port, A4(10) => 
                           X_Logic0_port, A4(9) => X_Logic0_port, A4(8) => 
                           X_Logic0_port, A4(7) => X_Logic0_port, A4(6) => 
                           X_Logic0_port, A4(5) => X_Logic0_port, A4(4) => 
                           X_Logic0_port, A4(3) => X_Logic0_port, A4(2) => 
                           X_Logic0_port, A4(1) => X_Logic0_port, A4(0) => 
                           X_Logic0_port, sel(2) => selVector_13_2_port, sel(1)
                           => selVector_13_1_port, sel(0) => 
                           selVector_13_0_port, O(63) => 
                           muxOutVector_13_63_port, O(62) => 
                           muxOutVector_13_62_port, O(61) => 
                           muxOutVector_13_61_port, O(60) => 
                           muxOutVector_13_60_port, O(59) => 
                           muxOutVector_13_59_port, O(58) => 
                           muxOutVector_13_58_port, O(57) => 
                           muxOutVector_13_57_port, O(56) => 
                           muxOutVector_13_56_port, O(55) => 
                           muxOutVector_13_55_port, O(54) => 
                           muxOutVector_13_54_port, O(53) => 
                           muxOutVector_13_53_port, O(52) => 
                           muxOutVector_13_52_port, O(51) => 
                           muxOutVector_13_51_port, O(50) => 
                           muxOutVector_13_50_port, O(49) => 
                           muxOutVector_13_49_port, O(48) => 
                           muxOutVector_13_48_port, O(47) => 
                           muxOutVector_13_47_port, O(46) => 
                           muxOutVector_13_46_port, O(45) => 
                           muxOutVector_13_45_port, O(44) => 
                           muxOutVector_13_44_port, O(43) => 
                           muxOutVector_13_43_port, O(42) => 
                           muxOutVector_13_42_port, O(41) => 
                           muxOutVector_13_41_port, O(40) => 
                           muxOutVector_13_40_port, O(39) => 
                           muxOutVector_13_39_port, O(38) => 
                           muxOutVector_13_38_port, O(37) => 
                           muxOutVector_13_37_port, O(36) => 
                           muxOutVector_13_36_port, O(35) => 
                           muxOutVector_13_35_port, O(34) => 
                           muxOutVector_13_34_port, O(33) => 
                           muxOutVector_13_33_port, O(32) => 
                           muxOutVector_13_32_port, O(31) => 
                           muxOutVector_13_31_port, O(30) => 
                           muxOutVector_13_30_port, O(29) => 
                           muxOutVector_13_29_port, O(28) => 
                           muxOutVector_13_28_port, O(27) => 
                           muxOutVector_13_27_port, O(26) => 
                           muxOutVector_13_26_port, O(25) => 
                           muxOutVector_13_25_port, O(24) => 
                           muxOutVector_13_24_port, O(23) => 
                           muxOutVector_13_23_port, O(22) => 
                           muxOutVector_13_22_port, O(21) => 
                           muxOutVector_13_21_port, O(20) => 
                           muxOutVector_13_20_port, O(19) => 
                           muxOutVector_13_19_port, O(18) => 
                           muxOutVector_13_18_port, O(17) => 
                           muxOutVector_13_17_port, O(16) => 
                           muxOutVector_13_16_port, O(15) => 
                           muxOutVector_13_15_port, O(14) => 
                           muxOutVector_13_14_port, O(13) => 
                           muxOutVector_13_13_port, O(12) => 
                           muxOutVector_13_12_port, O(11) => 
                           muxOutVector_13_11_port, O(10) => 
                           muxOutVector_13_10_port, O(9) => 
                           muxOutVector_13_9_port, O(8) => 
                           muxOutVector_13_8_port, O(7) => 
                           muxOutVector_13_7_port, O(6) => 
                           muxOutVector_13_6_port, O(5) => 
                           muxOutVector_13_5_port, O(4) => 
                           muxOutVector_13_4_port, O(3) => 
                           muxOutVector_13_3_port, O(2) => 
                           muxOutVector_13_2_port, O(1) => 
                           muxOutVector_13_1_port, O(0) => 
                           muxOutVector_13_0_port);
   eb_14 : BE_BLOCK_2 port map( b(2) => B(29), b(1) => B(28), b(0) => B(27), 
                           sel(2) => selVector_14_2_port, sel(1) => 
                           selVector_14_1_port, sel(0) => selVector_14_0_port);
   sum_14 : RCA_NBIT64_2 port map( A(63) => muxOutVector_14_63_port, A(62) => 
                           muxOutVector_14_62_port, A(61) => 
                           muxOutVector_14_61_port, A(60) => 
                           muxOutVector_14_60_port, A(59) => 
                           muxOutVector_14_59_port, A(58) => 
                           muxOutVector_14_58_port, A(57) => 
                           muxOutVector_14_57_port, A(56) => 
                           muxOutVector_14_56_port, A(55) => 
                           muxOutVector_14_55_port, A(54) => 
                           muxOutVector_14_54_port, A(53) => 
                           muxOutVector_14_53_port, A(52) => 
                           muxOutVector_14_52_port, A(51) => 
                           muxOutVector_14_51_port, A(50) => 
                           muxOutVector_14_50_port, A(49) => 
                           muxOutVector_14_49_port, A(48) => 
                           muxOutVector_14_48_port, A(47) => 
                           muxOutVector_14_47_port, A(46) => 
                           muxOutVector_14_46_port, A(45) => 
                           muxOutVector_14_45_port, A(44) => 
                           muxOutVector_14_44_port, A(43) => 
                           muxOutVector_14_43_port, A(42) => 
                           muxOutVector_14_42_port, A(41) => 
                           muxOutVector_14_41_port, A(40) => 
                           muxOutVector_14_40_port, A(39) => 
                           muxOutVector_14_39_port, A(38) => 
                           muxOutVector_14_38_port, A(37) => 
                           muxOutVector_14_37_port, A(36) => 
                           muxOutVector_14_36_port, A(35) => 
                           muxOutVector_14_35_port, A(34) => 
                           muxOutVector_14_34_port, A(33) => 
                           muxOutVector_14_33_port, A(32) => 
                           muxOutVector_14_32_port, A(31) => 
                           muxOutVector_14_31_port, A(30) => 
                           muxOutVector_14_30_port, A(29) => 
                           muxOutVector_14_29_port, A(28) => 
                           muxOutVector_14_28_port, A(27) => 
                           muxOutVector_14_27_port, A(26) => 
                           muxOutVector_14_26_port, A(25) => 
                           muxOutVector_14_25_port, A(24) => 
                           muxOutVector_14_24_port, A(23) => 
                           muxOutVector_14_23_port, A(22) => 
                           muxOutVector_14_22_port, A(21) => 
                           muxOutVector_14_21_port, A(20) => 
                           muxOutVector_14_20_port, A(19) => 
                           muxOutVector_14_19_port, A(18) => 
                           muxOutVector_14_18_port, A(17) => 
                           muxOutVector_14_17_port, A(16) => 
                           muxOutVector_14_16_port, A(15) => 
                           muxOutVector_14_15_port, A(14) => 
                           muxOutVector_14_14_port, A(13) => 
                           muxOutVector_14_13_port, A(12) => 
                           muxOutVector_14_12_port, A(11) => 
                           muxOutVector_14_11_port, A(10) => 
                           muxOutVector_14_10_port, A(9) => 
                           muxOutVector_14_9_port, A(8) => 
                           muxOutVector_14_8_port, A(7) => 
                           muxOutVector_14_7_port, A(6) => 
                           muxOutVector_14_6_port, A(5) => 
                           muxOutVector_14_5_port, A(4) => 
                           muxOutVector_14_4_port, A(3) => 
                           muxOutVector_14_3_port, A(2) => 
                           muxOutVector_14_2_port, A(1) => 
                           muxOutVector_14_1_port, A(0) => 
                           muxOutVector_14_0_port, B(63) => 
                           sumVector_13_63_port, B(62) => sumVector_13_62_port,
                           B(61) => sumVector_13_61_port, B(60) => 
                           sumVector_13_60_port, B(59) => sumVector_13_59_port,
                           B(58) => sumVector_13_58_port, B(57) => 
                           sumVector_13_57_port, B(56) => sumVector_13_56_port,
                           B(55) => sumVector_13_55_port, B(54) => 
                           sumVector_13_54_port, B(53) => sumVector_13_53_port,
                           B(52) => sumVector_13_52_port, B(51) => 
                           sumVector_13_51_port, B(50) => sumVector_13_50_port,
                           B(49) => sumVector_13_49_port, B(48) => 
                           sumVector_13_48_port, B(47) => sumVector_13_47_port,
                           B(46) => sumVector_13_46_port, B(45) => 
                           sumVector_13_45_port, B(44) => sumVector_13_44_port,
                           B(43) => sumVector_13_43_port, B(42) => 
                           sumVector_13_42_port, B(41) => sumVector_13_41_port,
                           B(40) => sumVector_13_40_port, B(39) => 
                           sumVector_13_39_port, B(38) => sumVector_13_38_port,
                           B(37) => sumVector_13_37_port, B(36) => 
                           sumVector_13_36_port, B(35) => sumVector_13_35_port,
                           B(34) => sumVector_13_34_port, B(33) => 
                           sumVector_13_33_port, B(32) => sumVector_13_32_port,
                           B(31) => sumVector_13_31_port, B(30) => 
                           sumVector_13_30_port, B(29) => sumVector_13_29_port,
                           B(28) => sumVector_13_28_port, B(27) => 
                           sumVector_13_27_port, B(26) => sumVector_13_26_port,
                           B(25) => sumVector_13_25_port, B(24) => 
                           sumVector_13_24_port, B(23) => sumVector_13_23_port,
                           B(22) => sumVector_13_22_port, B(21) => 
                           sumVector_13_21_port, B(20) => sumVector_13_20_port,
                           B(19) => sumVector_13_19_port, B(18) => 
                           sumVector_13_18_port, B(17) => sumVector_13_17_port,
                           B(16) => sumVector_13_16_port, B(15) => 
                           sumVector_13_15_port, B(14) => sumVector_13_14_port,
                           B(13) => sumVector_13_13_port, B(12) => 
                           sumVector_13_12_port, B(11) => sumVector_13_11_port,
                           B(10) => sumVector_13_10_port, B(9) => 
                           sumVector_13_9_port, B(8) => sumVector_13_8_port, 
                           B(7) => sumVector_13_7_port, B(6) => 
                           sumVector_13_6_port, B(5) => sumVector_13_5_port, 
                           B(4) => sumVector_13_4_port, B(3) => 
                           sumVector_13_3_port, B(2) => sumVector_13_2_port, 
                           B(1) => sumVector_13_1_port, B(0) => 
                           sumVector_13_0_port, Ci => X_Logic0_port, S(63) => 
                           sumVector_14_63_port, S(62) => sumVector_14_62_port,
                           S(61) => sumVector_14_61_port, S(60) => 
                           sumVector_14_60_port, S(59) => sumVector_14_59_port,
                           S(58) => sumVector_14_58_port, S(57) => 
                           sumVector_14_57_port, S(56) => sumVector_14_56_port,
                           S(55) => sumVector_14_55_port, S(54) => 
                           sumVector_14_54_port, S(53) => sumVector_14_53_port,
                           S(52) => sumVector_14_52_port, S(51) => 
                           sumVector_14_51_port, S(50) => sumVector_14_50_port,
                           S(49) => sumVector_14_49_port, S(48) => 
                           sumVector_14_48_port, S(47) => sumVector_14_47_port,
                           S(46) => sumVector_14_46_port, S(45) => 
                           sumVector_14_45_port, S(44) => sumVector_14_44_port,
                           S(43) => sumVector_14_43_port, S(42) => 
                           sumVector_14_42_port, S(41) => sumVector_14_41_port,
                           S(40) => sumVector_14_40_port, S(39) => 
                           sumVector_14_39_port, S(38) => sumVector_14_38_port,
                           S(37) => sumVector_14_37_port, S(36) => 
                           sumVector_14_36_port, S(35) => sumVector_14_35_port,
                           S(34) => sumVector_14_34_port, S(33) => 
                           sumVector_14_33_port, S(32) => sumVector_14_32_port,
                           S(31) => sumVector_14_31_port, S(30) => 
                           sumVector_14_30_port, S(29) => sumVector_14_29_port,
                           S(28) => sumVector_14_28_port, S(27) => 
                           sumVector_14_27_port, S(26) => sumVector_14_26_port,
                           S(25) => sumVector_14_25_port, S(24) => 
                           sumVector_14_24_port, S(23) => sumVector_14_23_port,
                           S(22) => sumVector_14_22_port, S(21) => 
                           sumVector_14_21_port, S(20) => sumVector_14_20_port,
                           S(19) => sumVector_14_19_port, S(18) => 
                           sumVector_14_18_port, S(17) => sumVector_14_17_port,
                           S(16) => sumVector_14_16_port, S(15) => 
                           sumVector_14_15_port, S(14) => sumVector_14_14_port,
                           S(13) => sumVector_14_13_port, S(12) => 
                           sumVector_14_12_port, S(11) => sumVector_14_11_port,
                           S(10) => sumVector_14_10_port, S(9) => 
                           sumVector_14_9_port, S(8) => sumVector_14_8_port, 
                           S(7) => sumVector_14_7_port, S(6) => 
                           sumVector_14_6_port, S(5) => sumVector_14_5_port, 
                           S(4) => sumVector_14_4_port, S(3) => 
                           sumVector_14_3_port, S(2) => sumVector_14_2_port, 
                           S(1) => sumVector_14_1_port, S(0) => 
                           sumVector_14_0_port, Co => n_1049);
   mux_14 : MUX_5TO1_NBIT64_2 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n123, A1(62) => n123, 
                           A1(61) => n123, A1(60) => n123, A1(59) => n123, 
                           A1(58) => n374, A1(57) => n367, A1(56) => n360, 
                           A1(55) => n353, A1(54) => n346, A1(53) => n339, 
                           A1(52) => n332, A1(51) => n325, A1(50) => n318, 
                           A1(49) => n311, A1(48) => n304, A1(47) => n297, 
                           A1(46) => n290, A1(45) => n283, A1(44) => n276, 
                           A1(43) => n269, A1(42) => n262, A1(41) => n255, 
                           A1(40) => n248, A1(39) => n241, A1(38) => n234, 
                           A1(37) => n227, A1(36) => n220, A1(35) => n213, 
                           A1(34) => n206, A1(33) => n199, A1(32) => n192, 
                           A1(31) => n186, A1(30) => n182, A1(29) => n176, 
                           A1(28) => A(0), A1(27) => X_Logic0_port, A1(26) => 
                           X_Logic0_port, A1(25) => X_Logic0_port, A1(24) => 
                           X_Logic0_port, A1(23) => X_Logic0_port, A1(22) => 
                           X_Logic0_port, A1(21) => X_Logic0_port, A1(20) => 
                           X_Logic0_port, A1(19) => X_Logic0_port, A1(18) => 
                           X_Logic0_port, A1(17) => X_Logic0_port, A1(16) => 
                           X_Logic0_port, A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(63) => n523, A2(62) => n523, 
                           A2(61) => n523, A2(60) => n523, A2(59) => n493, 
                           A2(58) => n489, A2(57) => n485, A2(56) => n481, 
                           A2(55) => n477, A2(54) => n473, A2(53) => n469, 
                           A2(52) => n465, A2(51) => n461, A2(50) => n457, 
                           A2(49) => n453, A2(48) => n449, A2(47) => n445, 
                           A2(46) => n441, A2(45) => n437, A2(44) => n433, 
                           A2(43) => n430, A2(42) => n426, A2(41) => n423, 
                           A2(40) => n420, A2(39) => n416, A2(38) => n412, 
                           A2(37) => n409, A2(36) => n405, A2(35) => n401, 
                           A2(34) => n398, A2(33) => n396, A2(32) => n392, 
                           A2(31) => n101, A2(30) => n387, A2(29) => n99, 
                           A2(28) => n168, A2(27) => X_Logic0_port, A2(26) => 
                           X_Logic0_port, A2(25) => X_Logic0_port, A2(24) => 
                           X_Logic0_port, A2(23) => X_Logic0_port, A2(22) => 
                           X_Logic0_port, A2(21) => X_Logic0_port, A2(20) => 
                           X_Logic0_port, A2(19) => X_Logic0_port, A2(18) => 
                           X_Logic0_port, A2(17) => X_Logic0_port, A2(16) => 
                           X_Logic0_port, A2(15) => X_Logic0_port, A2(14) => 
                           X_Logic0_port, A2(13) => X_Logic0_port, A2(12) => 
                           X_Logic0_port, A2(11) => X_Logic0_port, A2(10) => 
                           X_Logic0_port, A2(9) => X_Logic0_port, A2(8) => 
                           X_Logic0_port, A2(7) => X_Logic0_port, A2(6) => 
                           X_Logic0_port, A2(5) => X_Logic0_port, A2(4) => 
                           X_Logic0_port, A2(3) => X_Logic0_port, A2(2) => 
                           X_Logic0_port, A2(1) => X_Logic0_port, A2(0) => 
                           X_Logic0_port, A3(63) => n151, A3(62) => n151, 
                           A3(61) => n151, A3(60) => n151, A3(59) => n378, 
                           A3(58) => n371, A3(57) => n364, A3(56) => n357, 
                           A3(55) => n350, A3(54) => n343, A3(53) => n336, 
                           A3(52) => n329, A3(51) => n322, A3(50) => n315, 
                           A3(49) => n308, A3(48) => n301, A3(47) => n294, 
                           A3(46) => n287, A3(45) => n280, A3(44) => n273, 
                           A3(43) => n266, A3(42) => n259, A3(41) => n252, 
                           A3(40) => n245, A3(39) => n238, A3(38) => n231, 
                           A3(37) => n224, A3(36) => n217, A3(35) => n210, 
                           A3(34) => n203, A3(33) => n196, A3(32) => n186, 
                           A3(31) => n182, A3(30) => n176, A3(29) => A(0), 
                           A3(28) => X_Logic0_port, A3(27) => X_Logic0_port, 
                           A3(26) => X_Logic0_port, A3(25) => X_Logic0_port, 
                           A3(24) => X_Logic0_port, A3(23) => X_Logic0_port, 
                           A3(22) => X_Logic0_port, A3(21) => X_Logic0_port, 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n507, A4(62) => 
                           n507, A4(61) => n507, A4(60) => n492, A4(59) => n488
                           , A4(58) => n484, A4(57) => n480, A4(56) => n476, 
                           A4(55) => n472, A4(54) => n468, A4(53) => n464, 
                           A4(52) => n460, A4(51) => n456, A4(50) => n452, 
                           A4(49) => n448, A4(48) => n444, A4(47) => n440, 
                           A4(46) => n436, A4(45) => n432, A4(44) => n429, 
                           A4(43) => n425, A4(42) => n422, A4(41) => n419, 
                           A4(40) => n415, A4(39) => n411, A4(38) => n408, 
                           A4(37) => n404, A4(36) => n400, A4(35) => n105, 
                           A4(34) => n394, A4(33) => n391, A4(32) => n388, 
                           A4(31) => n386, A4(30) => n383, A4(29) => n167, 
                           A4(28) => X_Logic0_port, A4(27) => X_Logic0_port, 
                           A4(26) => X_Logic0_port, A4(25) => X_Logic0_port, 
                           A4(24) => X_Logic0_port, A4(23) => X_Logic0_port, 
                           A4(22) => X_Logic0_port, A4(21) => X_Logic0_port, 
                           A4(20) => X_Logic0_port, A4(19) => X_Logic0_port, 
                           A4(18) => X_Logic0_port, A4(17) => X_Logic0_port, 
                           A4(16) => X_Logic0_port, A4(15) => X_Logic0_port, 
                           A4(14) => X_Logic0_port, A4(13) => X_Logic0_port, 
                           A4(12) => X_Logic0_port, A4(11) => X_Logic0_port, 
                           A4(10) => X_Logic0_port, A4(9) => X_Logic0_port, 
                           A4(8) => X_Logic0_port, A4(7) => X_Logic0_port, 
                           A4(6) => X_Logic0_port, A4(5) => X_Logic0_port, 
                           A4(4) => X_Logic0_port, A4(3) => X_Logic0_port, 
                           A4(2) => X_Logic0_port, A4(1) => X_Logic0_port, 
                           A4(0) => X_Logic0_port, sel(2) => 
                           selVector_14_2_port, sel(1) => selVector_14_1_port, 
                           sel(0) => selVector_14_0_port, O(63) => 
                           muxOutVector_14_63_port, O(62) => 
                           muxOutVector_14_62_port, O(61) => 
                           muxOutVector_14_61_port, O(60) => 
                           muxOutVector_14_60_port, O(59) => 
                           muxOutVector_14_59_port, O(58) => 
                           muxOutVector_14_58_port, O(57) => 
                           muxOutVector_14_57_port, O(56) => 
                           muxOutVector_14_56_port, O(55) => 
                           muxOutVector_14_55_port, O(54) => 
                           muxOutVector_14_54_port, O(53) => 
                           muxOutVector_14_53_port, O(52) => 
                           muxOutVector_14_52_port, O(51) => 
                           muxOutVector_14_51_port, O(50) => 
                           muxOutVector_14_50_port, O(49) => 
                           muxOutVector_14_49_port, O(48) => 
                           muxOutVector_14_48_port, O(47) => 
                           muxOutVector_14_47_port, O(46) => 
                           muxOutVector_14_46_port, O(45) => 
                           muxOutVector_14_45_port, O(44) => 
                           muxOutVector_14_44_port, O(43) => 
                           muxOutVector_14_43_port, O(42) => 
                           muxOutVector_14_42_port, O(41) => 
                           muxOutVector_14_41_port, O(40) => 
                           muxOutVector_14_40_port, O(39) => 
                           muxOutVector_14_39_port, O(38) => 
                           muxOutVector_14_38_port, O(37) => 
                           muxOutVector_14_37_port, O(36) => 
                           muxOutVector_14_36_port, O(35) => 
                           muxOutVector_14_35_port, O(34) => 
                           muxOutVector_14_34_port, O(33) => 
                           muxOutVector_14_33_port, O(32) => 
                           muxOutVector_14_32_port, O(31) => 
                           muxOutVector_14_31_port, O(30) => 
                           muxOutVector_14_30_port, O(29) => 
                           muxOutVector_14_29_port, O(28) => 
                           muxOutVector_14_28_port, O(27) => 
                           muxOutVector_14_27_port, O(26) => 
                           muxOutVector_14_26_port, O(25) => 
                           muxOutVector_14_25_port, O(24) => 
                           muxOutVector_14_24_port, O(23) => 
                           muxOutVector_14_23_port, O(22) => 
                           muxOutVector_14_22_port, O(21) => 
                           muxOutVector_14_21_port, O(20) => 
                           muxOutVector_14_20_port, O(19) => 
                           muxOutVector_14_19_port, O(18) => 
                           muxOutVector_14_18_port, O(17) => 
                           muxOutVector_14_17_port, O(16) => 
                           muxOutVector_14_16_port, O(15) => 
                           muxOutVector_14_15_port, O(14) => 
                           muxOutVector_14_14_port, O(13) => 
                           muxOutVector_14_13_port, O(12) => 
                           muxOutVector_14_12_port, O(11) => 
                           muxOutVector_14_11_port, O(10) => 
                           muxOutVector_14_10_port, O(9) => 
                           muxOutVector_14_9_port, O(8) => 
                           muxOutVector_14_8_port, O(7) => 
                           muxOutVector_14_7_port, O(6) => 
                           muxOutVector_14_6_port, O(5) => 
                           muxOutVector_14_5_port, O(4) => 
                           muxOutVector_14_4_port, O(3) => 
                           muxOutVector_14_3_port, O(2) => 
                           muxOutVector_14_2_port, O(1) => 
                           muxOutVector_14_1_port, O(0) => 
                           muxOutVector_14_0_port);
   eb_15 : BE_BLOCK_1 port map( b(2) => B(31), b(1) => B(30), b(0) => B(29), 
                           sel(2) => selVector_15_2_port, sel(1) => 
                           selVector_15_1_port, sel(0) => selVector_15_0_port);
   sum_15 : RCA_NBIT64_1 port map( A(63) => muxOutVector_15_63_port, A(62) => 
                           muxOutVector_15_62_port, A(61) => 
                           muxOutVector_15_61_port, A(60) => 
                           muxOutVector_15_60_port, A(59) => 
                           muxOutVector_15_59_port, A(58) => 
                           muxOutVector_15_58_port, A(57) => 
                           muxOutVector_15_57_port, A(56) => 
                           muxOutVector_15_56_port, A(55) => 
                           muxOutVector_15_55_port, A(54) => 
                           muxOutVector_15_54_port, A(53) => 
                           muxOutVector_15_53_port, A(52) => 
                           muxOutVector_15_52_port, A(51) => 
                           muxOutVector_15_51_port, A(50) => 
                           muxOutVector_15_50_port, A(49) => 
                           muxOutVector_15_49_port, A(48) => 
                           muxOutVector_15_48_port, A(47) => 
                           muxOutVector_15_47_port, A(46) => 
                           muxOutVector_15_46_port, A(45) => 
                           muxOutVector_15_45_port, A(44) => 
                           muxOutVector_15_44_port, A(43) => 
                           muxOutVector_15_43_port, A(42) => 
                           muxOutVector_15_42_port, A(41) => 
                           muxOutVector_15_41_port, A(40) => 
                           muxOutVector_15_40_port, A(39) => 
                           muxOutVector_15_39_port, A(38) => 
                           muxOutVector_15_38_port, A(37) => 
                           muxOutVector_15_37_port, A(36) => 
                           muxOutVector_15_36_port, A(35) => 
                           muxOutVector_15_35_port, A(34) => 
                           muxOutVector_15_34_port, A(33) => 
                           muxOutVector_15_33_port, A(32) => 
                           muxOutVector_15_32_port, A(31) => 
                           muxOutVector_15_31_port, A(30) => 
                           muxOutVector_15_30_port, A(29) => 
                           muxOutVector_15_29_port, A(28) => 
                           muxOutVector_15_28_port, A(27) => 
                           muxOutVector_15_27_port, A(26) => 
                           muxOutVector_15_26_port, A(25) => 
                           muxOutVector_15_25_port, A(24) => 
                           muxOutVector_15_24_port, A(23) => 
                           muxOutVector_15_23_port, A(22) => 
                           muxOutVector_15_22_port, A(21) => 
                           muxOutVector_15_21_port, A(20) => 
                           muxOutVector_15_20_port, A(19) => 
                           muxOutVector_15_19_port, A(18) => 
                           muxOutVector_15_18_port, A(17) => 
                           muxOutVector_15_17_port, A(16) => 
                           muxOutVector_15_16_port, A(15) => 
                           muxOutVector_15_15_port, A(14) => 
                           muxOutVector_15_14_port, A(13) => 
                           muxOutVector_15_13_port, A(12) => 
                           muxOutVector_15_12_port, A(11) => 
                           muxOutVector_15_11_port, A(10) => 
                           muxOutVector_15_10_port, A(9) => 
                           muxOutVector_15_9_port, A(8) => 
                           muxOutVector_15_8_port, A(7) => 
                           muxOutVector_15_7_port, A(6) => 
                           muxOutVector_15_6_port, A(5) => 
                           muxOutVector_15_5_port, A(4) => 
                           muxOutVector_15_4_port, A(3) => 
                           muxOutVector_15_3_port, A(2) => 
                           muxOutVector_15_2_port, A(1) => 
                           muxOutVector_15_1_port, A(0) => 
                           muxOutVector_15_0_port, B(63) => 
                           sumVector_14_63_port, B(62) => sumVector_14_62_port,
                           B(61) => sumVector_14_61_port, B(60) => 
                           sumVector_14_60_port, B(59) => sumVector_14_59_port,
                           B(58) => sumVector_14_58_port, B(57) => 
                           sumVector_14_57_port, B(56) => sumVector_14_56_port,
                           B(55) => sumVector_14_55_port, B(54) => 
                           sumVector_14_54_port, B(53) => sumVector_14_53_port,
                           B(52) => sumVector_14_52_port, B(51) => 
                           sumVector_14_51_port, B(50) => sumVector_14_50_port,
                           B(49) => sumVector_14_49_port, B(48) => 
                           sumVector_14_48_port, B(47) => sumVector_14_47_port,
                           B(46) => sumVector_14_46_port, B(45) => 
                           sumVector_14_45_port, B(44) => sumVector_14_44_port,
                           B(43) => sumVector_14_43_port, B(42) => 
                           sumVector_14_42_port, B(41) => sumVector_14_41_port,
                           B(40) => sumVector_14_40_port, B(39) => 
                           sumVector_14_39_port, B(38) => sumVector_14_38_port,
                           B(37) => sumVector_14_37_port, B(36) => 
                           sumVector_14_36_port, B(35) => sumVector_14_35_port,
                           B(34) => sumVector_14_34_port, B(33) => 
                           sumVector_14_33_port, B(32) => sumVector_14_32_port,
                           B(31) => sumVector_14_31_port, B(30) => 
                           sumVector_14_30_port, B(29) => sumVector_14_29_port,
                           B(28) => sumVector_14_28_port, B(27) => 
                           sumVector_14_27_port, B(26) => sumVector_14_26_port,
                           B(25) => sumVector_14_25_port, B(24) => 
                           sumVector_14_24_port, B(23) => sumVector_14_23_port,
                           B(22) => sumVector_14_22_port, B(21) => 
                           sumVector_14_21_port, B(20) => sumVector_14_20_port,
                           B(19) => sumVector_14_19_port, B(18) => 
                           sumVector_14_18_port, B(17) => sumVector_14_17_port,
                           B(16) => sumVector_14_16_port, B(15) => 
                           sumVector_14_15_port, B(14) => sumVector_14_14_port,
                           B(13) => sumVector_14_13_port, B(12) => 
                           sumVector_14_12_port, B(11) => sumVector_14_11_port,
                           B(10) => sumVector_14_10_port, B(9) => 
                           sumVector_14_9_port, B(8) => sumVector_14_8_port, 
                           B(7) => sumVector_14_7_port, B(6) => 
                           sumVector_14_6_port, B(5) => sumVector_14_5_port, 
                           B(4) => sumVector_14_4_port, B(3) => 
                           sumVector_14_3_port, B(2) => sumVector_14_2_port, 
                           B(1) => sumVector_14_1_port, B(0) => 
                           sumVector_14_0_port, Ci => X_Logic0_port, S(63) => 
                           P(63), S(62) => P(62), S(61) => P(61), S(60) => 
                           P(60), S(59) => P(59), S(58) => P(58), S(57) => 
                           P(57), S(56) => P(56), S(55) => P(55), S(54) => 
                           P(54), S(53) => P(53), S(52) => P(52), S(51) => 
                           P(51), S(50) => P(50), S(49) => P(49), S(48) => 
                           P(48), S(47) => P(47), S(46) => P(46), S(45) => 
                           P(45), S(44) => P(44), S(43) => P(43), S(42) => 
                           P(42), S(41) => P(41), S(40) => P(40), S(39) => 
                           P(39), S(38) => P(38), S(37) => P(37), S(36) => 
                           P(36), S(35) => P(35), S(34) => P(34), S(33) => 
                           P(33), S(32) => P(32), S(31) => P(31), S(30) => 
                           P(30), S(29) => P(29), S(28) => P(28), S(27) => 
                           P(27), S(26) => P(26), S(25) => P(25), S(24) => 
                           P(24), S(23) => P(23), S(22) => P(22), S(21) => 
                           P(21), S(20) => P(20), S(19) => P(19), S(18) => 
                           P(18), S(17) => P(17), S(16) => P(16), S(15) => 
                           P(15), S(14) => P(14), S(13) => P(13), S(12) => 
                           P(12), S(11) => P(11), S(10) => P(10), S(9) => P(9),
                           S(8) => P(8), S(7) => P(7), S(6) => P(6), S(5) => 
                           P(5), S(4) => P(4), S(3) => P(3), S(2) => P(2), S(1)
                           => P(1), S(0) => P(0), Co => n_1050);
   mux_15 : MUX_5TO1_NBIT64_1 port map( A0(63) => X_Logic0_port, A0(62) => 
                           X_Logic0_port, A0(61) => X_Logic0_port, A0(60) => 
                           X_Logic0_port, A0(59) => X_Logic0_port, A0(58) => 
                           X_Logic0_port, A0(57) => X_Logic0_port, A0(56) => 
                           X_Logic0_port, A0(55) => X_Logic0_port, A0(54) => 
                           X_Logic0_port, A0(53) => X_Logic0_port, A0(52) => 
                           X_Logic0_port, A0(51) => X_Logic0_port, A0(50) => 
                           X_Logic0_port, A0(49) => X_Logic0_port, A0(48) => 
                           X_Logic0_port, A0(47) => X_Logic0_port, A0(46) => 
                           X_Logic0_port, A0(45) => X_Logic0_port, A0(44) => 
                           X_Logic0_port, A0(43) => X_Logic0_port, A0(42) => 
                           X_Logic0_port, A0(41) => X_Logic0_port, A0(40) => 
                           X_Logic0_port, A0(39) => X_Logic0_port, A0(38) => 
                           X_Logic0_port, A0(37) => X_Logic0_port, A0(36) => 
                           X_Logic0_port, A0(35) => X_Logic0_port, A0(34) => 
                           X_Logic0_port, A0(33) => X_Logic0_port, A0(32) => 
                           X_Logic0_port, A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(63) => n124, A1(62) => n124, 
                           A1(61) => n123, A1(60) => n376, A1(59) => n369, 
                           A1(58) => n362, A1(57) => n355, A1(56) => n348, 
                           A1(55) => n341, A1(54) => n334, A1(53) => n327, 
                           A1(52) => n320, A1(51) => n313, A1(50) => n306, 
                           A1(49) => n299, A1(48) => n292, A1(47) => n285, 
                           A1(46) => n278, A1(45) => n271, A1(44) => n264, 
                           A1(43) => n257, A1(42) => n250, A1(41) => n243, 
                           A1(40) => n236, A1(39) => n229, A1(38) => n222, 
                           A1(37) => n215, A1(36) => n208, A1(35) => n201, 
                           A1(34) => n194, A1(33) => n186, A1(32) => n182, 
                           A1(31) => n103, A1(30) => A(0), A1(29) => 
                           X_Logic0_port, A1(28) => X_Logic0_port, A1(27) => 
                           X_Logic0_port, A1(26) => X_Logic0_port, A1(25) => 
                           X_Logic0_port, A1(24) => X_Logic0_port, A1(23) => 
                           X_Logic0_port, A1(22) => X_Logic0_port, A1(21) => 
                           X_Logic0_port, A1(20) => X_Logic0_port, A1(19) => 
                           X_Logic0_port, A1(18) => X_Logic0_port, A1(17) => 
                           X_Logic0_port, A1(16) => X_Logic0_port, A1(15) => 
                           X_Logic0_port, A1(14) => X_Logic0_port, A1(13) => 
                           X_Logic0_port, A1(12) => X_Logic0_port, A1(11) => 
                           X_Logic0_port, A1(10) => X_Logic0_port, A1(9) => 
                           X_Logic0_port, A1(8) => X_Logic0_port, A1(7) => 
                           X_Logic0_port, A1(6) => X_Logic0_port, A1(5) => 
                           X_Logic0_port, A1(4) => X_Logic0_port, A1(3) => 
                           X_Logic0_port, A1(2) => X_Logic0_port, A1(1) => 
                           X_Logic0_port, A1(0) => X_Logic0_port, A2(63) => 
                           n524, A2(62) => n524, A2(61) => n493, A2(60) => n489
                           , A2(59) => n485, A2(58) => n481, A2(57) => n477, 
                           A2(56) => n473, A2(55) => n469, A2(54) => n465, 
                           A2(53) => n461, A2(52) => n457, A2(51) => n453, 
                           A2(50) => n449, A2(49) => n445, A2(48) => n441, 
                           A2(47) => n437, A2(46) => n433, A2(45) => n430, 
                           A2(44) => n426, A2(43) => n423, A2(42) => n420, 
                           A2(41) => n416, A2(40) => n412, A2(39) => n409, 
                           A2(38) => n405, A2(37) => n400, A2(36) => n104, 
                           A2(35) => n396, A2(34) => n392, A2(33) => n389, 
                           A2(32) => n387, A2(31) => n99, A2(30) => n168, 
                           A2(29) => X_Logic0_port, A2(28) => X_Logic0_port, 
                           A2(27) => X_Logic0_port, A2(26) => X_Logic0_port, 
                           A2(25) => X_Logic0_port, A2(24) => X_Logic0_port, 
                           A2(23) => X_Logic0_port, A2(22) => X_Logic0_port, 
                           A2(21) => X_Logic0_port, A2(20) => X_Logic0_port, 
                           A2(19) => X_Logic0_port, A2(18) => X_Logic0_port, 
                           A2(17) => X_Logic0_port, A2(16) => X_Logic0_port, 
                           A2(15) => X_Logic0_port, A2(14) => X_Logic0_port, 
                           A2(13) => X_Logic0_port, A2(12) => X_Logic0_port, 
                           A2(11) => X_Logic0_port, A2(10) => X_Logic0_port, 
                           A2(9) => X_Logic0_port, A2(8) => X_Logic0_port, 
                           A2(7) => X_Logic0_port, A2(6) => X_Logic0_port, 
                           A2(5) => X_Logic0_port, A2(4) => X_Logic0_port, 
                           A2(3) => X_Logic0_port, A2(2) => X_Logic0_port, 
                           A2(1) => X_Logic0_port, A2(0) => X_Logic0_port, 
                           A3(63) => n151, A3(62) => n151, A3(61) => n376, 
                           A3(60) => n369, A3(59) => n362, A3(58) => n355, 
                           A3(57) => n348, A3(56) => n341, A3(55) => n334, 
                           A3(54) => n327, A3(53) => n320, A3(52) => n313, 
                           A3(51) => n306, A3(50) => n299, A3(49) => n292, 
                           A3(48) => n285, A3(47) => n278, A3(46) => n271, 
                           A3(45) => n264, A3(44) => n257, A3(43) => n250, 
                           A3(42) => n243, A3(41) => n236, A3(40) => n229, 
                           A3(39) => n222, A3(38) => n215, A3(37) => n208, 
                           A3(36) => n201, A3(35) => n194, A3(34) => n186, 
                           A3(33) => n182, A3(32) => n176, A3(31) => A(0), 
                           A3(30) => X_Logic0_port, A3(29) => X_Logic0_port, 
                           A3(28) => X_Logic0_port, A3(27) => X_Logic0_port, 
                           A3(26) => X_Logic0_port, A3(25) => X_Logic0_port, 
                           A3(24) => X_Logic0_port, A3(23) => X_Logic0_port, 
                           A3(22) => X_Logic0_port, A3(21) => X_Logic0_port, 
                           A3(20) => X_Logic0_port, A3(19) => X_Logic0_port, 
                           A3(18) => X_Logic0_port, A3(17) => X_Logic0_port, 
                           A3(16) => X_Logic0_port, A3(15) => X_Logic0_port, 
                           A3(14) => X_Logic0_port, A3(13) => X_Logic0_port, 
                           A3(12) => X_Logic0_port, A3(11) => X_Logic0_port, 
                           A3(10) => X_Logic0_port, A3(9) => X_Logic0_port, 
                           A3(8) => X_Logic0_port, A3(7) => X_Logic0_port, 
                           A3(6) => X_Logic0_port, A3(5) => X_Logic0_port, 
                           A3(4) => X_Logic0_port, A3(3) => X_Logic0_port, 
                           A3(2) => X_Logic0_port, A3(1) => X_Logic0_port, 
                           A3(0) => X_Logic0_port, A4(63) => n507, A4(62) => 
                           n492, A4(61) => n488, A4(60) => n484, A4(59) => n480
                           , A4(58) => n476, A4(57) => n472, A4(56) => n468, 
                           A4(55) => n464, A4(54) => n460, A4(53) => n456, 
                           A4(52) => n452, A4(51) => n448, A4(50) => n444, 
                           A4(49) => n440, A4(48) => n436, A4(47) => n432, 
                           A4(46) => n429, A4(45) => n425, A4(44) => n422, 
                           A4(43) => n419, A4(42) => n415, A4(41) => n411, 
                           A4(40) => n408, A4(39) => n404, A4(38) => n400, 
                           A4(37) => n397, A4(36) => n396, A4(35) => n391, 
                           A4(34) => n100, A4(33) => n386, A4(32) => n385, 
                           A4(31) => n167, A4(30) => X_Logic0_port, A4(29) => 
                           X_Logic0_port, A4(28) => X_Logic0_port, A4(27) => 
                           X_Logic0_port, A4(26) => X_Logic0_port, A4(25) => 
                           X_Logic0_port, A4(24) => X_Logic0_port, A4(23) => 
                           X_Logic0_port, A4(22) => X_Logic0_port, A4(21) => 
                           X_Logic0_port, A4(20) => X_Logic0_port, A4(19) => 
                           X_Logic0_port, A4(18) => X_Logic0_port, A4(17) => 
                           X_Logic0_port, A4(16) => X_Logic0_port, A4(15) => 
                           X_Logic0_port, A4(14) => X_Logic0_port, A4(13) => 
                           X_Logic0_port, A4(12) => X_Logic0_port, A4(11) => 
                           X_Logic0_port, A4(10) => X_Logic0_port, A4(9) => 
                           X_Logic0_port, A4(8) => X_Logic0_port, A4(7) => 
                           X_Logic0_port, A4(6) => X_Logic0_port, A4(5) => 
                           X_Logic0_port, A4(4) => X_Logic0_port, A4(3) => 
                           X_Logic0_port, A4(2) => X_Logic0_port, A4(1) => 
                           X_Logic0_port, A4(0) => X_Logic0_port, sel(2) => 
                           selVector_15_2_port, sel(1) => selVector_15_1_port, 
                           sel(0) => selVector_15_0_port, O(63) => 
                           muxOutVector_15_63_port, O(62) => 
                           muxOutVector_15_62_port, O(61) => 
                           muxOutVector_15_61_port, O(60) => 
                           muxOutVector_15_60_port, O(59) => 
                           muxOutVector_15_59_port, O(58) => 
                           muxOutVector_15_58_port, O(57) => 
                           muxOutVector_15_57_port, O(56) => 
                           muxOutVector_15_56_port, O(55) => 
                           muxOutVector_15_55_port, O(54) => 
                           muxOutVector_15_54_port, O(53) => 
                           muxOutVector_15_53_port, O(52) => 
                           muxOutVector_15_52_port, O(51) => 
                           muxOutVector_15_51_port, O(50) => 
                           muxOutVector_15_50_port, O(49) => 
                           muxOutVector_15_49_port, O(48) => 
                           muxOutVector_15_48_port, O(47) => 
                           muxOutVector_15_47_port, O(46) => 
                           muxOutVector_15_46_port, O(45) => 
                           muxOutVector_15_45_port, O(44) => 
                           muxOutVector_15_44_port, O(43) => 
                           muxOutVector_15_43_port, O(42) => 
                           muxOutVector_15_42_port, O(41) => 
                           muxOutVector_15_41_port, O(40) => 
                           muxOutVector_15_40_port, O(39) => 
                           muxOutVector_15_39_port, O(38) => 
                           muxOutVector_15_38_port, O(37) => 
                           muxOutVector_15_37_port, O(36) => 
                           muxOutVector_15_36_port, O(35) => 
                           muxOutVector_15_35_port, O(34) => 
                           muxOutVector_15_34_port, O(33) => 
                           muxOutVector_15_33_port, O(32) => 
                           muxOutVector_15_32_port, O(31) => 
                           muxOutVector_15_31_port, O(30) => 
                           muxOutVector_15_30_port, O(29) => 
                           muxOutVector_15_29_port, O(28) => 
                           muxOutVector_15_28_port, O(27) => 
                           muxOutVector_15_27_port, O(26) => 
                           muxOutVector_15_26_port, O(25) => 
                           muxOutVector_15_25_port, O(24) => 
                           muxOutVector_15_24_port, O(23) => 
                           muxOutVector_15_23_port, O(22) => 
                           muxOutVector_15_22_port, O(21) => 
                           muxOutVector_15_21_port, O(20) => 
                           muxOutVector_15_20_port, O(19) => 
                           muxOutVector_15_19_port, O(18) => 
                           muxOutVector_15_18_port, O(17) => 
                           muxOutVector_15_17_port, O(16) => 
                           muxOutVector_15_16_port, O(15) => 
                           muxOutVector_15_15_port, O(14) => 
                           muxOutVector_15_14_port, O(13) => 
                           muxOutVector_15_13_port, O(12) => 
                           muxOutVector_15_12_port, O(11) => 
                           muxOutVector_15_11_port, O(10) => 
                           muxOutVector_15_10_port, O(9) => 
                           muxOutVector_15_9_port, O(8) => 
                           muxOutVector_15_8_port, O(7) => 
                           muxOutVector_15_7_port, O(6) => 
                           muxOutVector_15_6_port, O(5) => 
                           muxOutVector_15_5_port, O(4) => 
                           muxOutVector_15_4_port, O(3) => 
                           muxOutVector_15_3_port, O(2) => 
                           muxOutVector_15_2_port, O(1) => 
                           muxOutVector_15_1_port, O(0) => 
                           muxOutVector_15_0_port);
   r177 : BOOTHMUL_DW01_sub_0 port map( A(32) => n97, A(31) => n97, A(30) => 
                           n97, A(29) => n97, A(28) => n97, A(27) => n97, A(26)
                           => n97, A(25) => n97, A(24) => n97, A(23) => n97, 
                           A(22) => n97, A(21) => n97, A(20) => n97, A(19) => 
                           n97, A(18) => n97, A(17) => n97, A(16) => n97, A(15)
                           => n97, A(14) => n97, A(13) => n97, A(12) => n97, 
                           A(11) => n97, A(10) => n97, A(9) => n97, A(8) => n97
                           , A(7) => n97, A(6) => n97, A(5) => n97, A(4) => n97
                           , A(3) => n97, A(2) => n97, A(1) => n97, A(0) => n97
                           , B(32) => n381, B(31) => n557, B(30) => n374, B(29)
                           => n367, B(28) => n360, B(27) => n353, B(26) => n346
                           , B(25) => n339, B(24) => n332, B(23) => n325, B(22)
                           => n318, B(21) => n311, B(20) => n304, B(19) => n297
                           , B(18) => n290, B(17) => n283, B(16) => n276, B(15)
                           => n269, B(14) => n262, B(13) => n255, B(12) => n248
                           , B(11) => n241, B(10) => n234, B(9) => n227, B(8) 
                           => n220, B(7) => n213, B(6) => n206, B(5) => n199, 
                           B(4) => n192, B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n98, DIFF(32) => n3, 
                           DIFF(31) => n4, DIFF(30) => n5, DIFF(29) => n6, 
                           DIFF(28) => n7, DIFF(27) => n8, DIFF(26) => n9, 
                           DIFF(25) => n10, DIFF(24) => n11, DIFF(23) => n12, 
                           DIFF(22) => n13, DIFF(21) => n14, DIFF(20) => n15, 
                           DIFF(19) => n16, DIFF(18) => n17, DIFF(17) => n18, 
                           DIFF(16) => n19, DIFF(15) => n20, DIFF(14) => n21, 
                           DIFF(13) => n22, DIFF(12) => n23, DIFF(11) => n24, 
                           DIFF(10) => n25, DIFF(9) => n26, DIFF(8) => n27, 
                           DIFF(7) => n28, DIFF(6) => n29, DIFF(5) => n30, 
                           DIFF(4) => n31, DIFF(3) => n32, DIFF(2) => n33, 
                           DIFF(1) => n34, DIFF(0) => n35, CO => n_1051);
   U7 : BUF_X1 port map( A => A(2), Z => n178);
   U8 : BUF_X1 port map( A => A(17), Z => n283);
   U9 : BUF_X1 port map( A => A(18), Z => n290);
   U10 : BUF_X1 port map( A => A(19), Z => n297);
   U11 : BUF_X1 port map( A => A(20), Z => n304);
   U12 : BUF_X1 port map( A => n27, Z => n407);
   U13 : BUF_X1 port map( A => n25, Z => n414);
   U14 : BUF_X1 port map( A => n24, Z => n418);
   U15 : BUF_X1 port map( A => n21, Z => n428);
   U16 : BUF_X1 port map( A => n19, Z => n435);
   U17 : BUF_X1 port map( A => n18, Z => n439);
   U18 : BUF_X1 port map( A => n17, Z => n443);
   U19 : BUF_X1 port map( A => n16, Z => n447);
   U20 : BUF_X1 port map( A => n15, Z => n451);
   U21 : BUF_X1 port map( A => n14, Z => n455);
   U22 : BUF_X1 port map( A => n13, Z => n459);
   U23 : BUF_X1 port map( A => n12, Z => n463);
   U24 : BUF_X1 port map( A => n11, Z => n467);
   U25 : BUF_X1 port map( A => n10, Z => n471);
   U26 : BUF_X1 port map( A => n9, Z => n475);
   U27 : BUF_X1 port map( A => n8, Z => n479);
   U28 : BUF_X1 port map( A => n7, Z => n483);
   U29 : BUF_X1 port map( A => n6, Z => n487);
   U30 : BUF_X1 port map( A => n5, Z => n491);
   U31 : BUF_X1 port map( A => n4, Z => n495);
   U32 : BUF_X1 port map( A => n32, Z => n390);
   U33 : CLKBUF_X3 port map( A => n34, Z => n99);
   U34 : CLKBUF_X1 port map( A => n34, Z => n384);
   U35 : CLKBUF_X3 port map( A => n403, Z => n400);
   U36 : BUF_X2 port map( A => n403, Z => n401);
   U37 : BUF_X1 port map( A => n390, Z => n100);
   U38 : BUF_X1 port map( A => n390, Z => n101);
   U39 : BUF_X1 port map( A => n28, Z => n403);
   U40 : BUF_X1 port map( A => A(1), Z => n102);
   U41 : BUF_X2 port map( A => A(1), Z => n103);
   U42 : BUF_X2 port map( A => n399, Z => n105);
   U43 : BUF_X2 port map( A => A(1), Z => n176);
   U44 : BUF_X2 port map( A => n29, Z => n399);
   U45 : BUF_X1 port map( A => n399, Z => n104);
   U46 : BUF_X2 port map( A => n33, Z => n386);
   U47 : CLKBUF_X1 port map( A => n546, Z => n509);
   U48 : CLKBUF_X1 port map( A => n543, Z => n520);
   U49 : CLKBUF_X1 port map( A => n546, Z => n505);
   U50 : CLKBUF_X1 port map( A => n546, Z => n506);
   U51 : CLKBUF_X1 port map( A => n550, Z => n545);
   U52 : CLKBUF_X1 port map( A => n550, Z => n544);
   U53 : CLKBUF_X1 port map( A => n552, Z => n549);
   U54 : CLKBUF_X1 port map( A => n552, Z => n551);
   U55 : BUF_X2 port map( A => A(14), Z => n262);
   U56 : BUF_X1 port map( A => n550, Z => n543);
   U57 : BUF_X1 port map( A => n549, Z => n546);
   U58 : BUF_X1 port map( A => n551, Z => n540);
   U59 : BUF_X1 port map( A => n551, Z => n542);
   U60 : BUF_X1 port map( A => n551, Z => n541);
   U61 : BUF_X1 port map( A => n549, Z => n547);
   U62 : BUF_X1 port map( A => n552, Z => n550);
   U63 : CLKBUF_X1 port map( A => n495, Z => n494);
   U64 : CLKBUF_X1 port map( A => n31, Z => n393);
   U65 : BUF_X1 port map( A => n407, Z => n405);
   U66 : BUF_X2 port map( A => n26, Z => n409);
   U67 : CLKBUF_X1 port map( A => n399, Z => n398);
   U68 : CLKBUF_X1 port map( A => n26, Z => n410);
   U69 : CLKBUF_X1 port map( A => n23, Z => n421);
   U70 : CLKBUF_X1 port map( A => n22, Z => n424);
   U71 : CLKBUF_X1 port map( A => n439, Z => n438);
   U72 : BUF_X1 port map( A => n3, Z => n552);
   U73 : CLKBUF_X1 port map( A => n443, Z => n442);
   U74 : CLKBUF_X1 port map( A => n447, Z => n446);
   U75 : CLKBUF_X1 port map( A => n451, Z => n450);
   U76 : CLKBUF_X1 port map( A => n455, Z => n454);
   U77 : CLKBUF_X1 port map( A => n459, Z => n458);
   U78 : CLKBUF_X1 port map( A => n463, Z => n462);
   U79 : CLKBUF_X1 port map( A => n467, Z => n466);
   U80 : CLKBUF_X1 port map( A => n471, Z => n470);
   U81 : CLKBUF_X1 port map( A => n475, Z => n474);
   U82 : CLKBUF_X1 port map( A => n479, Z => n478);
   U83 : CLKBUF_X1 port map( A => n483, Z => n482);
   U84 : CLKBUF_X1 port map( A => n487, Z => n486);
   U85 : CLKBUF_X1 port map( A => n491, Z => n490);
   U86 : BUF_X1 port map( A => n382, Z => n117);
   U87 : BUF_X1 port map( A => n382, Z => n118);
   U88 : BUF_X1 port map( A => n382, Z => n119);
   U89 : BUF_X1 port map( A => n554, Z => n134);
   U90 : BUF_X1 port map( A => n556, Z => n166);
   U91 : BUF_X1 port map( A => n554, Z => n132);
   U92 : BUF_X1 port map( A => n555, Z => n147);
   U93 : BUF_X1 port map( A => n555, Z => n148);
   U94 : BUF_X1 port map( A => n553, Z => n382);
   U95 : BUF_X1 port map( A => n555, Z => n149);
   U96 : BUF_X1 port map( A => n554, Z => n133);
   U97 : BUF_X1 port map( A => n556, Z => n163);
   U98 : BUF_X1 port map( A => n556, Z => n164);
   U99 : BUF_X1 port map( A => n556, Z => n165);
   U100 : CLKBUF_X1 port map( A => n169, Z => n168);
   U101 : BUF_X1 port map( A => n559, Z => n554);
   U102 : BUF_X1 port map( A => n558, Z => n556);
   U103 : BUF_X1 port map( A => n558, Z => n555);
   U104 : BUF_X2 port map( A => A(7), Z => n213);
   U105 : BUF_X2 port map( A => A(8), Z => n220);
   U106 : BUF_X1 port map( A => A(12), Z => n248);
   U107 : BUF_X1 port map( A => A(13), Z => n255);
   U108 : BUF_X1 port map( A => A(15), Z => n269);
   U109 : BUF_X2 port map( A => A(16), Z => n276);
   U110 : BUF_X1 port map( A => A(21), Z => n311);
   U111 : BUF_X1 port map( A => A(22), Z => n318);
   U112 : BUF_X1 port map( A => A(23), Z => n325);
   U113 : BUF_X1 port map( A => A(24), Z => n332);
   U114 : BUF_X1 port map( A => A(25), Z => n339);
   U115 : BUF_X1 port map( A => A(26), Z => n346);
   U116 : BUF_X1 port map( A => A(27), Z => n353);
   U117 : BUF_X1 port map( A => A(28), Z => n360);
   U118 : BUF_X1 port map( A => A(29), Z => n367);
   U119 : BUF_X1 port map( A => A(30), Z => n374);
   U120 : BUF_X1 port map( A => A(31), Z => n559);
   U121 : BUF_X1 port map( A => A(31), Z => n558);
   U122 : BUF_X1 port map( A => n543, Z => n524);
   U123 : BUF_X1 port map( A => n546, Z => n507);
   U124 : BUF_X1 port map( A => n545, Z => n514);
   U125 : BUF_X1 port map( A => n544, Z => n515);
   U126 : BUF_X1 port map( A => n540, Z => n538);
   U127 : BUF_X1 port map( A => n545, Z => n511);
   U128 : BUF_X1 port map( A => n546, Z => n508);
   U129 : BUF_X1 port map( A => n542, Z => n525);
   U130 : BUF_X1 port map( A => n543, Z => n523);
   U131 : BUF_X1 port map( A => n543, Z => n522);
   U132 : BUF_X1 port map( A => n541, Z => n531);
   U133 : BUF_X1 port map( A => n545, Z => n512);
   U134 : BUF_X1 port map( A => n545, Z => n510);
   U135 : BUF_X1 port map( A => n541, Z => n530);
   U136 : BUF_X1 port map( A => n540, Z => n537);
   U137 : BUF_X1 port map( A => n542, Z => n528);
   U138 : BUF_X1 port map( A => n543, Z => n521);
   U139 : BUF_X1 port map( A => n544, Z => n517);
   U140 : BUF_X1 port map( A => n544, Z => n516);
   U141 : BUF_X1 port map( A => n540, Z => n536);
   U142 : BUF_X1 port map( A => n542, Z => n526);
   U143 : BUF_X1 port map( A => n548, Z => n497);
   U144 : BUF_X1 port map( A => n540, Z => n535);
   U145 : BUF_X1 port map( A => n547, Z => n503);
   U146 : BUF_X1 port map( A => n545, Z => n513);
   U147 : BUF_X1 port map( A => n548, Z => n496);
   U148 : BUF_X1 port map( A => n541, Z => n533);
   U149 : BUF_X1 port map( A => n548, Z => n499);
   U150 : BUF_X1 port map( A => n542, Z => n527);
   U151 : BUF_X1 port map( A => n548, Z => n498);
   U152 : BUF_X1 port map( A => n544, Z => n519);
   U153 : BUF_X1 port map( A => n542, Z => n529);
   U154 : BUF_X1 port map( A => n547, Z => n500);
   U155 : BUF_X1 port map( A => n541, Z => n532);
   U156 : BUF_X1 port map( A => n547, Z => n501);
   U157 : BUF_X1 port map( A => n544, Z => n518);
   U158 : BUF_X1 port map( A => n547, Z => n502);
   U159 : BUF_X1 port map( A => n541, Z => n534);
   U160 : BUF_X1 port map( A => n540, Z => n539);
   U161 : BUF_X1 port map( A => n547, Z => n504);
   U162 : BUF_X1 port map( A => n549, Z => n548);
   U163 : BUF_X1 port map( A => n393, Z => n391);
   U164 : BUF_X1 port map( A => n393, Z => n392);
   U165 : BUF_X1 port map( A => n495, Z => n493);
   U166 : BUF_X1 port map( A => n495, Z => n492);
   U167 : BUF_X1 port map( A => n117, Z => n114);
   U168 : BUF_X1 port map( A => n120, Z => n106);
   U169 : BUF_X1 port map( A => n118, Z => n113);
   U170 : BUF_X1 port map( A => n120, Z => n107);
   U171 : BUF_X1 port map( A => n119, Z => n108);
   U172 : BUF_X1 port map( A => n118, Z => n111);
   U173 : BUF_X1 port map( A => n119, Z => n109);
   U174 : BUF_X1 port map( A => n118, Z => n112);
   U175 : BUF_X1 port map( A => n117, Z => n116);
   U176 : BUF_X1 port map( A => n117, Z => n115);
   U177 : BUF_X1 port map( A => n119, Z => n110);
   U178 : BUF_X1 port map( A => n30, Z => n395);
   U179 : BUF_X1 port map( A => n418, Z => n416);
   U180 : BUF_X1 port map( A => n447, Z => n445);
   U181 : BUF_X2 port map( A => n390, Z => n389);
   U182 : BUF_X1 port map( A => n439, Z => n436);
   U183 : BUF_X1 port map( A => n23, Z => n420);
   U184 : BUF_X1 port map( A => n451, Z => n449);
   U185 : BUF_X1 port map( A => n443, Z => n440);
   U186 : BUF_X1 port map( A => n439, Z => n437);
   U187 : BUF_X1 port map( A => n399, Z => n397);
   U188 : BUF_X2 port map( A => n30, Z => n394);
   U189 : BUF_X1 port map( A => n22, Z => n423);
   U190 : BUF_X1 port map( A => n455, Z => n453);
   U191 : BUF_X1 port map( A => n20, Z => n429);
   U192 : BUF_X1 port map( A => n447, Z => n444);
   U193 : BUF_X1 port map( A => n414, Z => n412);
   U194 : BUF_X1 port map( A => n443, Z => n441);
   U195 : BUF_X1 port map( A => n20, Z => n430);
   U196 : BUF_X1 port map( A => n428, Z => n426);
   U197 : CLKBUF_X1 port map( A => n418, Z => n415);
   U198 : BUF_X1 port map( A => n459, Z => n457);
   U199 : BUF_X1 port map( A => n451, Z => n448);
   U200 : BUF_X1 port map( A => n23, Z => n419);
   U201 : BUF_X1 port map( A => n407, Z => n404);
   U202 : BUF_X1 port map( A => n463, Z => n461);
   U203 : BUF_X1 port map( A => n455, Z => n452);
   U204 : BUF_X1 port map( A => n435, Z => n433);
   U205 : BUF_X1 port map( A => n22, Z => n422);
   U206 : BUF_X1 port map( A => n26, Z => n408);
   U207 : BUF_X1 port map( A => n467, Z => n465);
   U208 : BUF_X1 port map( A => n459, Z => n456);
   U209 : CLKBUF_X1 port map( A => n428, Z => n425);
   U210 : BUF_X1 port map( A => n471, Z => n469);
   U211 : CLKBUF_X1 port map( A => n414, Z => n411);
   U212 : BUF_X1 port map( A => n463, Z => n460);
   U213 : BUF_X1 port map( A => n475, Z => n473);
   U214 : CLKBUF_X1 port map( A => n435, Z => n432);
   U215 : BUF_X1 port map( A => n467, Z => n464);
   U216 : BUF_X1 port map( A => n479, Z => n477);
   U217 : CLKBUF_X1 port map( A => n403, Z => n402);
   U218 : BUF_X1 port map( A => n471, Z => n468);
   U219 : BUF_X1 port map( A => n483, Z => n481);
   U220 : CLKBUF_X1 port map( A => n407, Z => n406);
   U221 : BUF_X1 port map( A => n475, Z => n472);
   U222 : BUF_X1 port map( A => n487, Z => n485);
   U223 : BUF_X1 port map( A => n479, Z => n476);
   U224 : BUF_X1 port map( A => n491, Z => n489);
   U225 : BUF_X1 port map( A => n483, Z => n480);
   U226 : BUF_X1 port map( A => n20, Z => n431);
   U227 : CLKBUF_X1 port map( A => n418, Z => n417);
   U228 : BUF_X1 port map( A => n487, Z => n484);
   U229 : BUF_X1 port map( A => n491, Z => n488);
   U230 : CLKBUF_X1 port map( A => n414, Z => n413);
   U231 : CLKBUF_X1 port map( A => n428, Z => n427);
   U232 : CLKBUF_X1 port map( A => n435, Z => n434);
   U233 : BUF_X1 port map( A => n134, Z => n124);
   U234 : BUF_X1 port map( A => n166, Z => n151);
   U235 : BUF_X1 port map( A => n132, Z => n130);
   U236 : BUF_X1 port map( A => n147, Z => n146);
   U237 : BUF_X1 port map( A => n148, Z => n142);
   U238 : BUF_X1 port map( A => n150, Z => n137);
   U239 : BUF_X1 port map( A => n149, Z => n140);
   U240 : BUF_X1 port map( A => n147, Z => n145);
   U241 : BUF_X1 port map( A => n382, Z => n120);
   U242 : BUF_X1 port map( A => n149, Z => n138);
   U243 : BUF_X1 port map( A => n134, Z => n125);
   U244 : BUF_X1 port map( A => n148, Z => n143);
   U245 : BUF_X1 port map( A => n149, Z => n139);
   U246 : BUF_X1 port map( A => n132, Z => n131);
   U247 : BUF_X1 port map( A => n147, Z => n144);
   U248 : BUF_X1 port map( A => n133, Z => n127);
   U249 : BUF_X1 port map( A => n133, Z => n128);
   U250 : BUF_X1 port map( A => n163, Z => n162);
   U251 : BUF_X1 port map( A => n133, Z => n126);
   U252 : BUF_X1 port map( A => n135, Z => n121);
   U253 : BUF_X1 port map( A => n163, Z => n160);
   U254 : BUF_X1 port map( A => n163, Z => n161);
   U255 : BUF_X1 port map( A => n148, Z => n141);
   U256 : BUF_X1 port map( A => n132, Z => n129);
   U257 : BUF_X1 port map( A => n164, Z => n158);
   U258 : BUF_X1 port map( A => n164, Z => n159);
   U259 : BUF_X1 port map( A => n164, Z => n157);
   U260 : BUF_X1 port map( A => n165, Z => n156);
   U261 : BUF_X1 port map( A => n135, Z => n122);
   U262 : BUF_X1 port map( A => n165, Z => n155);
   U263 : BUF_X1 port map( A => n150, Z => n136);
   U264 : BUF_X1 port map( A => n165, Z => n154);
   U265 : BUF_X1 port map( A => n166, Z => n153);
   U266 : BUF_X1 port map( A => n166, Z => n152);
   U267 : BUF_X1 port map( A => n134, Z => n123);
   U268 : BUF_X1 port map( A => n553, Z => n381);
   U269 : BUF_X1 port map( A => n555, Z => n150);
   U270 : BUF_X1 port map( A => n554, Z => n135);
   U271 : BUF_X1 port map( A => n34, Z => n383);
   U272 : CLKBUF_X1 port map( A => n34, Z => n385);
   U273 : BUF_X1 port map( A => n169, Z => n167);
   U274 : BUF_X1 port map( A => n559, Z => n553);
   U275 : BUF_X1 port map( A => n558, Z => n557);
   U276 : BUF_X1 port map( A => A(6), Z => n206);
   U277 : BUF_X2 port map( A => A(11), Z => n241);
   U278 : BUF_X1 port map( A => A(4), Z => n195);
   U279 : BUF_X1 port map( A => A(4), Z => n192);
   U280 : BUF_X1 port map( A => A(5), Z => n199);
   U281 : BUF_X1 port map( A => A(1), Z => n177);
   U282 : BUF_X1 port map( A => A(4), Z => n197);
   U283 : BUF_X1 port map( A => A(1), Z => n174);
   U284 : BUF_X1 port map( A => A(9), Z => n227);
   U285 : BUF_X1 port map( A => A(10), Z => n234);
   U286 : BUF_X1 port map( A => A(5), Z => n204);
   U287 : BUF_X1 port map( A => A(7), Z => n216);
   U288 : BUF_X1 port map( A => A(5), Z => n202);
   U289 : BUF_X1 port map( A => A(8), Z => n223);
   U290 : BUF_X1 port map( A => A(6), Z => n211);
   U291 : BUF_X1 port map( A => A(6), Z => n209);
   U292 : BUF_X1 port map( A => A(7), Z => n218);
   U293 : BUF_X1 port map( A => A(9), Z => n230);
   U294 : BUF_X1 port map( A => A(4), Z => n196);
   U295 : BUF_X1 port map( A => A(8), Z => n225);
   U296 : BUF_X1 port map( A => A(10), Z => n237);
   U297 : BUF_X1 port map( A => n35, Z => n169);
   U298 : BUF_X1 port map( A => A(5), Z => n203);
   U299 : BUF_X1 port map( A => A(9), Z => n232);
   U300 : BUF_X1 port map( A => A(11), Z => n244);
   U301 : BUF_X1 port map( A => A(6), Z => n210);
   U302 : BUF_X1 port map( A => A(10), Z => n239);
   U303 : BUF_X1 port map( A => A(12), Z => n251);
   U304 : BUF_X1 port map( A => A(11), Z => n246);
   U305 : BUF_X1 port map( A => A(7), Z => n217);
   U306 : BUF_X1 port map( A => A(13), Z => n258);
   U307 : BUF_X1 port map( A => A(1), Z => n175);
   U308 : BUF_X1 port map( A => A(8), Z => n224);
   U309 : BUF_X1 port map( A => A(12), Z => n253);
   U310 : BUF_X1 port map( A => A(14), Z => n265);
   U311 : BUF_X1 port map( A => A(4), Z => n193);
   U312 : BUF_X1 port map( A => A(9), Z => n231);
   U313 : BUF_X1 port map( A => A(13), Z => n260);
   U314 : BUF_X1 port map( A => A(15), Z => n272);
   U315 : BUF_X1 port map( A => A(5), Z => n200);
   U316 : BUF_X1 port map( A => A(10), Z => n238);
   U317 : BUF_X1 port map( A => A(14), Z => n267);
   U318 : BUF_X1 port map( A => A(16), Z => n279);
   U319 : BUF_X1 port map( A => A(6), Z => n207);
   U320 : BUF_X1 port map( A => A(11), Z => n245);
   U321 : BUF_X1 port map( A => A(15), Z => n274);
   U322 : BUF_X1 port map( A => A(17), Z => n286);
   U323 : BUF_X1 port map( A => A(7), Z => n214);
   U324 : BUF_X1 port map( A => A(12), Z => n252);
   U325 : BUF_X1 port map( A => A(16), Z => n281);
   U326 : BUF_X1 port map( A => A(18), Z => n293);
   U327 : BUF_X1 port map( A => A(8), Z => n221);
   U328 : BUF_X1 port map( A => A(13), Z => n259);
   U329 : BUF_X1 port map( A => A(17), Z => n288);
   U330 : BUF_X1 port map( A => A(19), Z => n300);
   U331 : BUF_X1 port map( A => A(9), Z => n228);
   U332 : BUF_X1 port map( A => A(14), Z => n266);
   U333 : BUF_X1 port map( A => A(18), Z => n295);
   U334 : BUF_X1 port map( A => A(20), Z => n307);
   U335 : BUF_X1 port map( A => A(10), Z => n235);
   U336 : BUF_X1 port map( A => A(15), Z => n273);
   U337 : BUF_X1 port map( A => A(19), Z => n302);
   U338 : BUF_X1 port map( A => A(21), Z => n314);
   U339 : BUF_X1 port map( A => A(11), Z => n242);
   U340 : BUF_X1 port map( A => A(16), Z => n280);
   U341 : BUF_X1 port map( A => A(20), Z => n309);
   U342 : BUF_X1 port map( A => A(2), Z => n182);
   U343 : BUF_X1 port map( A => A(22), Z => n321);
   U344 : BUF_X1 port map( A => A(4), Z => n194);
   U345 : BUF_X1 port map( A => A(3), Z => n186);
   U346 : BUF_X1 port map( A => A(12), Z => n249);
   U347 : BUF_X1 port map( A => A(17), Z => n287);
   U348 : BUF_X1 port map( A => A(21), Z => n316);
   U349 : BUF_X1 port map( A => A(23), Z => n328);
   U350 : BUF_X1 port map( A => A(5), Z => n201);
   U351 : BUF_X1 port map( A => A(13), Z => n256);
   U352 : BUF_X1 port map( A => A(24), Z => n335);
   U353 : BUF_X1 port map( A => A(22), Z => n323);
   U354 : BUF_X1 port map( A => A(18), Z => n294);
   U355 : BUF_X1 port map( A => A(6), Z => n208);
   U356 : BUF_X1 port map( A => A(14), Z => n263);
   U357 : BUF_X1 port map( A => A(19), Z => n301);
   U358 : BUF_X1 port map( A => A(23), Z => n330);
   U359 : BUF_X1 port map( A => A(25), Z => n342);
   U360 : BUF_X1 port map( A => A(7), Z => n215);
   U361 : BUF_X1 port map( A => A(4), Z => n198);
   U362 : BUF_X1 port map( A => A(15), Z => n270);
   U363 : BUF_X1 port map( A => A(20), Z => n308);
   U364 : BUF_X1 port map( A => A(24), Z => n337);
   U365 : BUF_X1 port map( A => A(26), Z => n349);
   U366 : BUF_X1 port map( A => A(8), Z => n222);
   U367 : BUF_X1 port map( A => A(5), Z => n205);
   U368 : BUF_X1 port map( A => A(16), Z => n277);
   U369 : BUF_X1 port map( A => A(21), Z => n315);
   U370 : BUF_X1 port map( A => A(25), Z => n344);
   U371 : BUF_X1 port map( A => A(27), Z => n356);
   U372 : BUF_X1 port map( A => A(9), Z => n229);
   U373 : BUF_X1 port map( A => A(6), Z => n212);
   U374 : BUF_X1 port map( A => A(17), Z => n284);
   U375 : BUF_X1 port map( A => A(26), Z => n351);
   U376 : BUF_X1 port map( A => A(22), Z => n322);
   U377 : BUF_X1 port map( A => A(28), Z => n363);
   U378 : BUF_X1 port map( A => A(10), Z => n236);
   U379 : BUF_X1 port map( A => A(7), Z => n219);
   U380 : BUF_X1 port map( A => A(18), Z => n291);
   U381 : BUF_X1 port map( A => A(23), Z => n329);
   U382 : BUF_X1 port map( A => A(27), Z => n358);
   U383 : BUF_X1 port map( A => A(29), Z => n370);
   U384 : BUF_X1 port map( A => A(11), Z => n243);
   U385 : BUF_X1 port map( A => A(8), Z => n226);
   U386 : BUF_X1 port map( A => A(19), Z => n298);
   U387 : BUF_X1 port map( A => A(28), Z => n364);
   U388 : BUF_X1 port map( A => A(24), Z => n336);
   U389 : BUF_X1 port map( A => A(28), Z => n365);
   U390 : BUF_X1 port map( A => A(30), Z => n377);
   U391 : BUF_X1 port map( A => A(12), Z => n250);
   U392 : BUF_X1 port map( A => A(9), Z => n233);
   U393 : BUF_X1 port map( A => A(20), Z => n305);
   U394 : BUF_X1 port map( A => A(29), Z => n372);
   U395 : BUF_X1 port map( A => A(25), Z => n343);
   U396 : BUF_X1 port map( A => A(13), Z => n257);
   U397 : BUF_X1 port map( A => A(10), Z => n240);
   U398 : BUF_X1 port map( A => A(21), Z => n312);
   U399 : BUF_X1 port map( A => A(26), Z => n350);
   U400 : BUF_X1 port map( A => A(30), Z => n379);
   U401 : BUF_X1 port map( A => A(14), Z => n264);
   U402 : BUF_X1 port map( A => A(11), Z => n247);
   U403 : BUF_X1 port map( A => A(22), Z => n319);
   U404 : BUF_X1 port map( A => A(27), Z => n357);
   U405 : BUF_X1 port map( A => A(15), Z => n271);
   U406 : BUF_X1 port map( A => A(12), Z => n254);
   U407 : BUF_X1 port map( A => A(23), Z => n326);
   U408 : BUF_X1 port map( A => A(16), Z => n278);
   U409 : BUF_X1 port map( A => A(13), Z => n261);
   U410 : BUF_X1 port map( A => A(24), Z => n333);
   U411 : BUF_X1 port map( A => A(29), Z => n371);
   U412 : BUF_X1 port map( A => A(17), Z => n285);
   U413 : BUF_X1 port map( A => A(14), Z => n268);
   U414 : BUF_X1 port map( A => A(25), Z => n340);
   U415 : BUF_X1 port map( A => A(30), Z => n378);
   U416 : BUF_X1 port map( A => A(18), Z => n292);
   U417 : BUF_X1 port map( A => A(15), Z => n275);
   U418 : BUF_X1 port map( A => A(26), Z => n347);
   U419 : BUF_X1 port map( A => A(19), Z => n299);
   U420 : BUF_X1 port map( A => A(16), Z => n282);
   U421 : BUF_X1 port map( A => A(27), Z => n354);
   U422 : BUF_X1 port map( A => A(20), Z => n306);
   U423 : BUF_X1 port map( A => A(17), Z => n289);
   U424 : BUF_X1 port map( A => A(28), Z => n361);
   U425 : BUF_X1 port map( A => A(21), Z => n313);
   U426 : BUF_X1 port map( A => A(18), Z => n296);
   U427 : BUF_X1 port map( A => A(29), Z => n368);
   U428 : BUF_X1 port map( A => A(22), Z => n320);
   U429 : BUF_X1 port map( A => A(19), Z => n303);
   U430 : BUF_X1 port map( A => A(30), Z => n375);
   U431 : BUF_X1 port map( A => A(23), Z => n327);
   U432 : BUF_X1 port map( A => A(20), Z => n310);
   U433 : BUF_X1 port map( A => A(24), Z => n334);
   U434 : BUF_X1 port map( A => A(21), Z => n317);
   U435 : BUF_X1 port map( A => A(25), Z => n341);
   U436 : BUF_X1 port map( A => A(22), Z => n324);
   U437 : BUF_X1 port map( A => A(26), Z => n348);
   U438 : BUF_X1 port map( A => A(23), Z => n331);
   U439 : BUF_X1 port map( A => A(27), Z => n355);
   U440 : BUF_X1 port map( A => A(24), Z => n338);
   U441 : BUF_X1 port map( A => A(28), Z => n362);
   U442 : BUF_X1 port map( A => A(25), Z => n345);
   U443 : BUF_X1 port map( A => A(29), Z => n369);
   U444 : BUF_X1 port map( A => A(26), Z => n352);
   U445 : BUF_X1 port map( A => A(30), Z => n376);
   U446 : BUF_X1 port map( A => A(27), Z => n359);
   U447 : BUF_X1 port map( A => A(28), Z => n366);
   U448 : BUF_X1 port map( A => A(29), Z => n373);
   U449 : BUF_X1 port map( A => A(30), Z => n380);
   U450 : BUF_X1 port map( A => A(3), Z => n170);
   U451 : BUF_X1 port map( A => A(3), Z => n171);
   U452 : BUF_X1 port map( A => A(3), Z => n185);
   U453 : BUF_X1 port map( A => A(3), Z => n190);
   U454 : BUF_X1 port map( A => A(3), Z => n188);
   U455 : BUF_X1 port map( A => A(3), Z => n191);
   U456 : BUF_X1 port map( A => A(3), Z => n187);
   U457 : BUF_X1 port map( A => A(3), Z => n189);
   U458 : BUF_X1 port map( A => A(2), Z => n172);
   U459 : BUF_X1 port map( A => A(2), Z => n173);
   U460 : BUF_X1 port map( A => A(2), Z => n184);
   U461 : BUF_X1 port map( A => A(2), Z => n183);
   U462 : BUF_X1 port map( A => A(2), Z => n181);
   U463 : BUF_X1 port map( A => A(2), Z => n180);
   U464 : BUF_X1 port map( A => A(2), Z => n179);
   U465 : BUF_X2 port map( A => n33, Z => n387);
   U466 : BUF_X1 port map( A => n390, Z => n388);
   U467 : BUF_X2 port map( A => n30, Z => n396);

end SYN_MIXED;

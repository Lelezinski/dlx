LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.constants.ALL;

ENTITY CARRY_GENERATOR IS
	-- Generics changed to NBIT_PER_BLOCK and NBLOCKS to match the other TBs. 
	GENERIC (
		NBIT_PER_BLOCK : INTEGER := CARRY_SELECT_NBIT;
		NBLOCKS : INTEGER := SUM_GENERATOR_NBLOCK);
	PORT (
		A : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
		Cin : IN STD_LOGIC;
		Co : OUT STD_LOGIC_VECTOR(NBLOCKS - 1 DOWNTO 0));
END CARRY_GENERATOR;

ARCHITECTURE STRUCTURAL OF CARRY_GENERATOR IS
-- Structural description of the Carry Generator Block

	-- Top PG Network
	COMPONENT PG_NETWORK IS
		GENERIC (
			NBIT_PER_BLOCK : INTEGER := CARRY_SELECT_NBIT;
			NBLOCKS : INTEGER := SUM_GENERATOR_NBLOCK);
		PORT (
			A : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
			Cin : IN STD_LOGIC;
			g : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS DOWNTO 0);
			p : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS DOWNTO 0));
	END COMPONENT;

	-- G Block: General GENERATE
	COMPONENT G_BLOCK IS
		PORT (
			G_left : IN STD_LOGIC;
			P_left : IN STD_LOGIC;
			G_right : IN STD_LOGIC;

			G_out : OUT STD_LOGIC);
	END COMPONENT;

	-- PG Block: General PROPAGATE and General GENERATE
	COMPONENT PG_BLOCK IS
		PORT (
			G_left : IN STD_LOGIC;
			P_left : IN STD_LOGIC;
			G_right : IN STD_LOGIC;
			P_right : IN STD_LOGIC;

			P_out : OUT STD_LOGIC;
			G_out : OUT STD_LOGIC);
	END COMPONENT;	

	-- Arrays
		-- TODO: WRITE arrays

BEGIN
-- Components Istantiation
	pgn: PG_NETWORK
	GENERIC MAP(CARRY_SELECT_NBIT, SUM_GENERATOR_NBLOCK)
	PORT MAP(A, B, Cin, , ); -- TODO: FIX

	-- TODO: WRITE generate...

END STRUCTURAL;
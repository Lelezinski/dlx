
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file;

architecture SYN_A of register_file is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal NEXT_REGISTERS_0_63_port, NEXT_REGISTERS_0_62_port, 
      NEXT_REGISTERS_0_61_port, NEXT_REGISTERS_0_60_port, 
      NEXT_REGISTERS_0_59_port, NEXT_REGISTERS_0_58_port, 
      NEXT_REGISTERS_0_57_port, NEXT_REGISTERS_0_56_port, 
      NEXT_REGISTERS_0_55_port, NEXT_REGISTERS_0_54_port, 
      NEXT_REGISTERS_0_53_port, NEXT_REGISTERS_0_52_port, 
      NEXT_REGISTERS_0_51_port, NEXT_REGISTERS_0_50_port, 
      NEXT_REGISTERS_0_49_port, NEXT_REGISTERS_0_48_port, 
      NEXT_REGISTERS_0_47_port, NEXT_REGISTERS_0_46_port, 
      NEXT_REGISTERS_0_45_port, NEXT_REGISTERS_0_44_port, 
      NEXT_REGISTERS_0_43_port, NEXT_REGISTERS_0_42_port, 
      NEXT_REGISTERS_0_41_port, NEXT_REGISTERS_0_40_port, 
      NEXT_REGISTERS_0_39_port, NEXT_REGISTERS_0_38_port, 
      NEXT_REGISTERS_0_37_port, NEXT_REGISTERS_0_36_port, 
      NEXT_REGISTERS_0_35_port, NEXT_REGISTERS_0_34_port, 
      NEXT_REGISTERS_0_33_port, NEXT_REGISTERS_0_32_port, 
      NEXT_REGISTERS_0_31_port, NEXT_REGISTERS_0_30_port, 
      NEXT_REGISTERS_0_29_port, NEXT_REGISTERS_0_28_port, 
      NEXT_REGISTERS_0_27_port, NEXT_REGISTERS_0_26_port, 
      NEXT_REGISTERS_0_25_port, NEXT_REGISTERS_0_24_port, 
      NEXT_REGISTERS_0_23_port, NEXT_REGISTERS_0_22_port, 
      NEXT_REGISTERS_0_21_port, NEXT_REGISTERS_0_20_port, 
      NEXT_REGISTERS_0_19_port, NEXT_REGISTERS_0_18_port, 
      NEXT_REGISTERS_0_17_port, NEXT_REGISTERS_0_16_port, 
      NEXT_REGISTERS_0_15_port, NEXT_REGISTERS_0_14_port, 
      NEXT_REGISTERS_0_13_port, NEXT_REGISTERS_0_12_port, 
      NEXT_REGISTERS_0_11_port, NEXT_REGISTERS_0_10_port, 
      NEXT_REGISTERS_0_9_port, NEXT_REGISTERS_0_8_port, NEXT_REGISTERS_0_7_port
      , NEXT_REGISTERS_0_6_port, NEXT_REGISTERS_0_5_port, 
      NEXT_REGISTERS_0_4_port, NEXT_REGISTERS_0_3_port, NEXT_REGISTERS_0_2_port
      , NEXT_REGISTERS_0_1_port, NEXT_REGISTERS_0_0_port, 
      NEXT_REGISTERS_1_63_port, NEXT_REGISTERS_1_62_port, 
      NEXT_REGISTERS_1_61_port, NEXT_REGISTERS_1_60_port, 
      NEXT_REGISTERS_1_59_port, NEXT_REGISTERS_1_58_port, 
      NEXT_REGISTERS_1_57_port, NEXT_REGISTERS_1_56_port, 
      NEXT_REGISTERS_1_55_port, NEXT_REGISTERS_1_54_port, 
      NEXT_REGISTERS_1_53_port, NEXT_REGISTERS_1_52_port, 
      NEXT_REGISTERS_1_51_port, NEXT_REGISTERS_1_50_port, 
      NEXT_REGISTERS_1_49_port, NEXT_REGISTERS_1_48_port, 
      NEXT_REGISTERS_1_47_port, NEXT_REGISTERS_1_46_port, 
      NEXT_REGISTERS_1_45_port, NEXT_REGISTERS_1_44_port, 
      NEXT_REGISTERS_1_43_port, NEXT_REGISTERS_1_42_port, 
      NEXT_REGISTERS_1_41_port, NEXT_REGISTERS_1_40_port, 
      NEXT_REGISTERS_1_39_port, NEXT_REGISTERS_1_38_port, 
      NEXT_REGISTERS_1_37_port, NEXT_REGISTERS_1_36_port, 
      NEXT_REGISTERS_1_35_port, NEXT_REGISTERS_1_34_port, 
      NEXT_REGISTERS_1_33_port, NEXT_REGISTERS_1_32_port, 
      NEXT_REGISTERS_1_31_port, NEXT_REGISTERS_1_30_port, 
      NEXT_REGISTERS_1_29_port, NEXT_REGISTERS_1_28_port, 
      NEXT_REGISTERS_1_27_port, NEXT_REGISTERS_1_26_port, 
      NEXT_REGISTERS_1_25_port, NEXT_REGISTERS_1_24_port, 
      NEXT_REGISTERS_1_23_port, NEXT_REGISTERS_1_22_port, 
      NEXT_REGISTERS_1_21_port, NEXT_REGISTERS_1_20_port, 
      NEXT_REGISTERS_1_19_port, NEXT_REGISTERS_1_18_port, 
      NEXT_REGISTERS_1_17_port, NEXT_REGISTERS_1_16_port, 
      NEXT_REGISTERS_1_15_port, NEXT_REGISTERS_1_14_port, 
      NEXT_REGISTERS_1_13_port, NEXT_REGISTERS_1_12_port, 
      NEXT_REGISTERS_1_11_port, NEXT_REGISTERS_1_10_port, 
      NEXT_REGISTERS_1_9_port, NEXT_REGISTERS_1_8_port, NEXT_REGISTERS_1_7_port
      , NEXT_REGISTERS_1_6_port, NEXT_REGISTERS_1_5_port, 
      NEXT_REGISTERS_1_4_port, NEXT_REGISTERS_1_3_port, NEXT_REGISTERS_1_2_port
      , NEXT_REGISTERS_1_1_port, NEXT_REGISTERS_1_0_port, 
      NEXT_REGISTERS_2_63_port, NEXT_REGISTERS_2_62_port, 
      NEXT_REGISTERS_2_61_port, NEXT_REGISTERS_2_60_port, 
      NEXT_REGISTERS_2_59_port, NEXT_REGISTERS_2_58_port, 
      NEXT_REGISTERS_2_57_port, NEXT_REGISTERS_2_56_port, 
      NEXT_REGISTERS_2_55_port, NEXT_REGISTERS_2_54_port, 
      NEXT_REGISTERS_2_53_port, NEXT_REGISTERS_2_52_port, 
      NEXT_REGISTERS_2_51_port, NEXT_REGISTERS_2_50_port, 
      NEXT_REGISTERS_2_49_port, NEXT_REGISTERS_2_48_port, 
      NEXT_REGISTERS_2_47_port, NEXT_REGISTERS_2_46_port, 
      NEXT_REGISTERS_2_45_port, NEXT_REGISTERS_2_44_port, 
      NEXT_REGISTERS_2_43_port, NEXT_REGISTERS_2_42_port, 
      NEXT_REGISTERS_2_41_port, NEXT_REGISTERS_2_40_port, 
      NEXT_REGISTERS_2_39_port, NEXT_REGISTERS_2_38_port, 
      NEXT_REGISTERS_2_37_port, NEXT_REGISTERS_2_36_port, 
      NEXT_REGISTERS_2_35_port, NEXT_REGISTERS_2_34_port, 
      NEXT_REGISTERS_2_33_port, NEXT_REGISTERS_2_32_port, 
      NEXT_REGISTERS_2_31_port, NEXT_REGISTERS_2_30_port, 
      NEXT_REGISTERS_2_29_port, NEXT_REGISTERS_2_28_port, 
      NEXT_REGISTERS_2_27_port, NEXT_REGISTERS_2_26_port, 
      NEXT_REGISTERS_2_25_port, NEXT_REGISTERS_2_24_port, 
      NEXT_REGISTERS_2_23_port, NEXT_REGISTERS_2_22_port, 
      NEXT_REGISTERS_2_21_port, NEXT_REGISTERS_2_20_port, 
      NEXT_REGISTERS_2_19_port, NEXT_REGISTERS_2_18_port, 
      NEXT_REGISTERS_2_17_port, NEXT_REGISTERS_2_16_port, 
      NEXT_REGISTERS_2_15_port, NEXT_REGISTERS_2_14_port, 
      NEXT_REGISTERS_2_13_port, NEXT_REGISTERS_2_12_port, 
      NEXT_REGISTERS_2_11_port, NEXT_REGISTERS_2_10_port, 
      NEXT_REGISTERS_2_9_port, NEXT_REGISTERS_2_8_port, NEXT_REGISTERS_2_7_port
      , NEXT_REGISTERS_2_6_port, NEXT_REGISTERS_2_5_port, 
      NEXT_REGISTERS_2_4_port, NEXT_REGISTERS_2_3_port, NEXT_REGISTERS_2_2_port
      , NEXT_REGISTERS_2_1_port, NEXT_REGISTERS_2_0_port, 
      NEXT_REGISTERS_3_63_port, NEXT_REGISTERS_3_62_port, 
      NEXT_REGISTERS_3_61_port, NEXT_REGISTERS_3_60_port, 
      NEXT_REGISTERS_3_59_port, NEXT_REGISTERS_3_58_port, 
      NEXT_REGISTERS_3_57_port, NEXT_REGISTERS_3_56_port, 
      NEXT_REGISTERS_3_55_port, NEXT_REGISTERS_3_54_port, 
      NEXT_REGISTERS_3_53_port, NEXT_REGISTERS_3_52_port, 
      NEXT_REGISTERS_3_51_port, NEXT_REGISTERS_3_50_port, 
      NEXT_REGISTERS_3_49_port, NEXT_REGISTERS_3_48_port, 
      NEXT_REGISTERS_3_47_port, NEXT_REGISTERS_3_46_port, 
      NEXT_REGISTERS_3_45_port, NEXT_REGISTERS_3_44_port, 
      NEXT_REGISTERS_3_43_port, NEXT_REGISTERS_3_42_port, 
      NEXT_REGISTERS_3_41_port, NEXT_REGISTERS_3_40_port, 
      NEXT_REGISTERS_3_39_port, NEXT_REGISTERS_3_38_port, 
      NEXT_REGISTERS_3_37_port, NEXT_REGISTERS_3_36_port, 
      NEXT_REGISTERS_3_35_port, NEXT_REGISTERS_3_34_port, 
      NEXT_REGISTERS_3_33_port, NEXT_REGISTERS_3_32_port, 
      NEXT_REGISTERS_3_31_port, NEXT_REGISTERS_3_30_port, 
      NEXT_REGISTERS_3_29_port, NEXT_REGISTERS_3_28_port, 
      NEXT_REGISTERS_3_27_port, NEXT_REGISTERS_3_26_port, 
      NEXT_REGISTERS_3_25_port, NEXT_REGISTERS_3_24_port, 
      NEXT_REGISTERS_3_23_port, NEXT_REGISTERS_3_22_port, 
      NEXT_REGISTERS_3_21_port, NEXT_REGISTERS_3_20_port, 
      NEXT_REGISTERS_3_19_port, NEXT_REGISTERS_3_18_port, 
      NEXT_REGISTERS_3_17_port, NEXT_REGISTERS_3_16_port, 
      NEXT_REGISTERS_3_15_port, NEXT_REGISTERS_3_14_port, 
      NEXT_REGISTERS_3_13_port, NEXT_REGISTERS_3_12_port, 
      NEXT_REGISTERS_3_11_port, NEXT_REGISTERS_3_10_port, 
      NEXT_REGISTERS_3_9_port, NEXT_REGISTERS_3_8_port, NEXT_REGISTERS_3_7_port
      , NEXT_REGISTERS_3_6_port, NEXT_REGISTERS_3_5_port, 
      NEXT_REGISTERS_3_4_port, NEXT_REGISTERS_3_3_port, NEXT_REGISTERS_3_2_port
      , NEXT_REGISTERS_3_1_port, NEXT_REGISTERS_3_0_port, 
      NEXT_REGISTERS_4_63_port, NEXT_REGISTERS_4_62_port, 
      NEXT_REGISTERS_4_61_port, NEXT_REGISTERS_4_60_port, 
      NEXT_REGISTERS_4_59_port, NEXT_REGISTERS_4_58_port, 
      NEXT_REGISTERS_4_57_port, NEXT_REGISTERS_4_56_port, 
      NEXT_REGISTERS_4_55_port, NEXT_REGISTERS_4_54_port, 
      NEXT_REGISTERS_4_53_port, NEXT_REGISTERS_4_52_port, 
      NEXT_REGISTERS_4_51_port, NEXT_REGISTERS_4_50_port, 
      NEXT_REGISTERS_4_49_port, NEXT_REGISTERS_4_48_port, 
      NEXT_REGISTERS_4_47_port, NEXT_REGISTERS_4_46_port, 
      NEXT_REGISTERS_4_45_port, NEXT_REGISTERS_4_44_port, 
      NEXT_REGISTERS_4_43_port, NEXT_REGISTERS_4_42_port, 
      NEXT_REGISTERS_4_41_port, NEXT_REGISTERS_4_40_port, 
      NEXT_REGISTERS_4_39_port, NEXT_REGISTERS_4_38_port, 
      NEXT_REGISTERS_4_37_port, NEXT_REGISTERS_4_36_port, 
      NEXT_REGISTERS_4_35_port, NEXT_REGISTERS_4_34_port, 
      NEXT_REGISTERS_4_33_port, NEXT_REGISTERS_4_32_port, 
      NEXT_REGISTERS_4_31_port, NEXT_REGISTERS_4_30_port, 
      NEXT_REGISTERS_4_29_port, NEXT_REGISTERS_4_28_port, 
      NEXT_REGISTERS_4_27_port, NEXT_REGISTERS_4_26_port, 
      NEXT_REGISTERS_4_25_port, NEXT_REGISTERS_4_24_port, 
      NEXT_REGISTERS_4_23_port, NEXT_REGISTERS_4_22_port, 
      NEXT_REGISTERS_4_21_port, NEXT_REGISTERS_4_20_port, 
      NEXT_REGISTERS_4_19_port, NEXT_REGISTERS_4_18_port, 
      NEXT_REGISTERS_4_17_port, NEXT_REGISTERS_4_16_port, 
      NEXT_REGISTERS_4_15_port, NEXT_REGISTERS_4_14_port, 
      NEXT_REGISTERS_4_13_port, NEXT_REGISTERS_4_12_port, 
      NEXT_REGISTERS_4_11_port, NEXT_REGISTERS_4_10_port, 
      NEXT_REGISTERS_4_9_port, NEXT_REGISTERS_4_8_port, NEXT_REGISTERS_4_7_port
      , NEXT_REGISTERS_4_6_port, NEXT_REGISTERS_4_5_port, 
      NEXT_REGISTERS_4_4_port, NEXT_REGISTERS_4_3_port, NEXT_REGISTERS_4_2_port
      , NEXT_REGISTERS_4_1_port, NEXT_REGISTERS_4_0_port, 
      NEXT_REGISTERS_5_63_port, NEXT_REGISTERS_5_62_port, 
      NEXT_REGISTERS_5_61_port, NEXT_REGISTERS_5_60_port, 
      NEXT_REGISTERS_5_59_port, NEXT_REGISTERS_5_58_port, 
      NEXT_REGISTERS_5_57_port, NEXT_REGISTERS_5_56_port, 
      NEXT_REGISTERS_5_55_port, NEXT_REGISTERS_5_54_port, 
      NEXT_REGISTERS_5_53_port, NEXT_REGISTERS_5_52_port, 
      NEXT_REGISTERS_5_51_port, NEXT_REGISTERS_5_50_port, 
      NEXT_REGISTERS_5_49_port, NEXT_REGISTERS_5_48_port, 
      NEXT_REGISTERS_5_47_port, NEXT_REGISTERS_5_46_port, 
      NEXT_REGISTERS_5_45_port, NEXT_REGISTERS_5_44_port, 
      NEXT_REGISTERS_5_43_port, NEXT_REGISTERS_5_42_port, 
      NEXT_REGISTERS_5_41_port, NEXT_REGISTERS_5_40_port, 
      NEXT_REGISTERS_5_39_port, NEXT_REGISTERS_5_38_port, 
      NEXT_REGISTERS_5_37_port, NEXT_REGISTERS_5_36_port, 
      NEXT_REGISTERS_5_35_port, NEXT_REGISTERS_5_34_port, 
      NEXT_REGISTERS_5_33_port, NEXT_REGISTERS_5_32_port, 
      NEXT_REGISTERS_5_31_port, NEXT_REGISTERS_5_30_port, 
      NEXT_REGISTERS_5_29_port, NEXT_REGISTERS_5_28_port, 
      NEXT_REGISTERS_5_27_port, NEXT_REGISTERS_5_26_port, 
      NEXT_REGISTERS_5_25_port, NEXT_REGISTERS_5_24_port, 
      NEXT_REGISTERS_5_23_port, NEXT_REGISTERS_5_22_port, 
      NEXT_REGISTERS_5_21_port, NEXT_REGISTERS_5_20_port, 
      NEXT_REGISTERS_5_19_port, NEXT_REGISTERS_5_18_port, 
      NEXT_REGISTERS_5_17_port, NEXT_REGISTERS_5_16_port, 
      NEXT_REGISTERS_5_15_port, NEXT_REGISTERS_5_14_port, 
      NEXT_REGISTERS_5_13_port, NEXT_REGISTERS_5_12_port, 
      NEXT_REGISTERS_5_11_port, NEXT_REGISTERS_5_10_port, 
      NEXT_REGISTERS_5_9_port, NEXT_REGISTERS_5_8_port, NEXT_REGISTERS_5_7_port
      , NEXT_REGISTERS_5_6_port, NEXT_REGISTERS_5_5_port, 
      NEXT_REGISTERS_5_4_port, NEXT_REGISTERS_5_3_port, NEXT_REGISTERS_5_2_port
      , NEXT_REGISTERS_5_1_port, NEXT_REGISTERS_5_0_port, 
      NEXT_REGISTERS_6_63_port, NEXT_REGISTERS_6_62_port, 
      NEXT_REGISTERS_6_61_port, NEXT_REGISTERS_6_60_port, 
      NEXT_REGISTERS_6_59_port, NEXT_REGISTERS_6_58_port, 
      NEXT_REGISTERS_6_57_port, NEXT_REGISTERS_6_56_port, 
      NEXT_REGISTERS_6_55_port, NEXT_REGISTERS_6_54_port, 
      NEXT_REGISTERS_6_53_port, NEXT_REGISTERS_6_52_port, 
      NEXT_REGISTERS_6_51_port, NEXT_REGISTERS_6_50_port, 
      NEXT_REGISTERS_6_49_port, NEXT_REGISTERS_6_48_port, 
      NEXT_REGISTERS_6_47_port, NEXT_REGISTERS_6_46_port, 
      NEXT_REGISTERS_6_45_port, NEXT_REGISTERS_6_44_port, 
      NEXT_REGISTERS_6_43_port, NEXT_REGISTERS_6_42_port, 
      NEXT_REGISTERS_6_41_port, NEXT_REGISTERS_6_40_port, 
      NEXT_REGISTERS_6_39_port, NEXT_REGISTERS_6_38_port, 
      NEXT_REGISTERS_6_37_port, NEXT_REGISTERS_6_36_port, 
      NEXT_REGISTERS_6_35_port, NEXT_REGISTERS_6_34_port, 
      NEXT_REGISTERS_6_33_port, NEXT_REGISTERS_6_32_port, 
      NEXT_REGISTERS_6_31_port, NEXT_REGISTERS_6_30_port, 
      NEXT_REGISTERS_6_29_port, NEXT_REGISTERS_6_28_port, 
      NEXT_REGISTERS_6_27_port, NEXT_REGISTERS_6_26_port, 
      NEXT_REGISTERS_6_25_port, NEXT_REGISTERS_6_24_port, 
      NEXT_REGISTERS_6_23_port, NEXT_REGISTERS_6_22_port, 
      NEXT_REGISTERS_6_21_port, NEXT_REGISTERS_6_20_port, 
      NEXT_REGISTERS_6_19_port, NEXT_REGISTERS_6_18_port, 
      NEXT_REGISTERS_6_17_port, NEXT_REGISTERS_6_16_port, 
      NEXT_REGISTERS_6_15_port, NEXT_REGISTERS_6_14_port, 
      NEXT_REGISTERS_6_13_port, NEXT_REGISTERS_6_12_port, 
      NEXT_REGISTERS_6_11_port, NEXT_REGISTERS_6_10_port, 
      NEXT_REGISTERS_6_9_port, NEXT_REGISTERS_6_8_port, NEXT_REGISTERS_6_7_port
      , NEXT_REGISTERS_6_6_port, NEXT_REGISTERS_6_5_port, 
      NEXT_REGISTERS_6_4_port, NEXT_REGISTERS_6_3_port, NEXT_REGISTERS_6_2_port
      , NEXT_REGISTERS_6_1_port, NEXT_REGISTERS_6_0_port, 
      NEXT_REGISTERS_7_63_port, NEXT_REGISTERS_7_62_port, 
      NEXT_REGISTERS_7_61_port, NEXT_REGISTERS_7_60_port, 
      NEXT_REGISTERS_7_59_port, NEXT_REGISTERS_7_58_port, 
      NEXT_REGISTERS_7_57_port, NEXT_REGISTERS_7_56_port, 
      NEXT_REGISTERS_7_55_port, NEXT_REGISTERS_7_54_port, 
      NEXT_REGISTERS_7_53_port, NEXT_REGISTERS_7_52_port, 
      NEXT_REGISTERS_7_51_port, NEXT_REGISTERS_7_50_port, 
      NEXT_REGISTERS_7_49_port, NEXT_REGISTERS_7_48_port, 
      NEXT_REGISTERS_7_47_port, NEXT_REGISTERS_7_46_port, 
      NEXT_REGISTERS_7_45_port, NEXT_REGISTERS_7_44_port, 
      NEXT_REGISTERS_7_43_port, NEXT_REGISTERS_7_42_port, 
      NEXT_REGISTERS_7_41_port, NEXT_REGISTERS_7_40_port, 
      NEXT_REGISTERS_7_39_port, NEXT_REGISTERS_7_38_port, 
      NEXT_REGISTERS_7_37_port, NEXT_REGISTERS_7_36_port, 
      NEXT_REGISTERS_7_35_port, NEXT_REGISTERS_7_34_port, 
      NEXT_REGISTERS_7_33_port, NEXT_REGISTERS_7_32_port, 
      NEXT_REGISTERS_7_31_port, NEXT_REGISTERS_7_30_port, 
      NEXT_REGISTERS_7_29_port, NEXT_REGISTERS_7_28_port, 
      NEXT_REGISTERS_7_27_port, NEXT_REGISTERS_7_26_port, 
      NEXT_REGISTERS_7_25_port, NEXT_REGISTERS_7_24_port, 
      NEXT_REGISTERS_7_23_port, NEXT_REGISTERS_7_22_port, 
      NEXT_REGISTERS_7_21_port, NEXT_REGISTERS_7_20_port, 
      NEXT_REGISTERS_7_19_port, NEXT_REGISTERS_7_18_port, 
      NEXT_REGISTERS_7_17_port, NEXT_REGISTERS_7_16_port, 
      NEXT_REGISTERS_7_15_port, NEXT_REGISTERS_7_14_port, 
      NEXT_REGISTERS_7_13_port, NEXT_REGISTERS_7_12_port, 
      NEXT_REGISTERS_7_11_port, NEXT_REGISTERS_7_10_port, 
      NEXT_REGISTERS_7_9_port, NEXT_REGISTERS_7_8_port, NEXT_REGISTERS_7_7_port
      , NEXT_REGISTERS_7_6_port, NEXT_REGISTERS_7_5_port, 
      NEXT_REGISTERS_7_4_port, NEXT_REGISTERS_7_3_port, NEXT_REGISTERS_7_2_port
      , NEXT_REGISTERS_7_1_port, NEXT_REGISTERS_7_0_port, 
      NEXT_REGISTERS_8_63_port, NEXT_REGISTERS_8_62_port, 
      NEXT_REGISTERS_8_61_port, NEXT_REGISTERS_8_60_port, 
      NEXT_REGISTERS_8_59_port, NEXT_REGISTERS_8_58_port, 
      NEXT_REGISTERS_8_57_port, NEXT_REGISTERS_8_56_port, 
      NEXT_REGISTERS_8_55_port, NEXT_REGISTERS_8_54_port, 
      NEXT_REGISTERS_8_53_port, NEXT_REGISTERS_8_52_port, 
      NEXT_REGISTERS_8_51_port, NEXT_REGISTERS_8_50_port, 
      NEXT_REGISTERS_8_49_port, NEXT_REGISTERS_8_48_port, 
      NEXT_REGISTERS_8_47_port, NEXT_REGISTERS_8_46_port, 
      NEXT_REGISTERS_8_45_port, NEXT_REGISTERS_8_44_port, 
      NEXT_REGISTERS_8_43_port, NEXT_REGISTERS_8_42_port, 
      NEXT_REGISTERS_8_41_port, NEXT_REGISTERS_8_40_port, 
      NEXT_REGISTERS_8_39_port, NEXT_REGISTERS_8_38_port, 
      NEXT_REGISTERS_8_37_port, NEXT_REGISTERS_8_36_port, 
      NEXT_REGISTERS_8_35_port, NEXT_REGISTERS_8_34_port, 
      NEXT_REGISTERS_8_33_port, NEXT_REGISTERS_8_32_port, 
      NEXT_REGISTERS_8_31_port, NEXT_REGISTERS_8_30_port, 
      NEXT_REGISTERS_8_29_port, NEXT_REGISTERS_8_28_port, 
      NEXT_REGISTERS_8_27_port, NEXT_REGISTERS_8_26_port, 
      NEXT_REGISTERS_8_25_port, NEXT_REGISTERS_8_24_port, 
      NEXT_REGISTERS_8_23_port, NEXT_REGISTERS_8_22_port, 
      NEXT_REGISTERS_8_21_port, NEXT_REGISTERS_8_20_port, 
      NEXT_REGISTERS_8_19_port, NEXT_REGISTERS_8_18_port, 
      NEXT_REGISTERS_8_17_port, NEXT_REGISTERS_8_16_port, 
      NEXT_REGISTERS_8_15_port, NEXT_REGISTERS_8_14_port, 
      NEXT_REGISTERS_8_13_port, NEXT_REGISTERS_8_12_port, 
      NEXT_REGISTERS_8_11_port, NEXT_REGISTERS_8_10_port, 
      NEXT_REGISTERS_8_9_port, NEXT_REGISTERS_8_8_port, NEXT_REGISTERS_8_7_port
      , NEXT_REGISTERS_8_6_port, NEXT_REGISTERS_8_5_port, 
      NEXT_REGISTERS_8_4_port, NEXT_REGISTERS_8_3_port, NEXT_REGISTERS_8_2_port
      , NEXT_REGISTERS_8_1_port, NEXT_REGISTERS_8_0_port, 
      NEXT_REGISTERS_9_63_port, NEXT_REGISTERS_9_62_port, 
      NEXT_REGISTERS_9_61_port, NEXT_REGISTERS_9_60_port, 
      NEXT_REGISTERS_9_59_port, NEXT_REGISTERS_9_58_port, 
      NEXT_REGISTERS_9_57_port, NEXT_REGISTERS_9_56_port, 
      NEXT_REGISTERS_9_55_port, NEXT_REGISTERS_9_54_port, 
      NEXT_REGISTERS_9_53_port, NEXT_REGISTERS_9_52_port, 
      NEXT_REGISTERS_9_51_port, NEXT_REGISTERS_9_50_port, 
      NEXT_REGISTERS_9_49_port, NEXT_REGISTERS_9_48_port, 
      NEXT_REGISTERS_9_47_port, NEXT_REGISTERS_9_46_port, 
      NEXT_REGISTERS_9_45_port, NEXT_REGISTERS_9_44_port, 
      NEXT_REGISTERS_9_43_port, NEXT_REGISTERS_9_42_port, 
      NEXT_REGISTERS_9_41_port, NEXT_REGISTERS_9_40_port, 
      NEXT_REGISTERS_9_39_port, NEXT_REGISTERS_9_38_port, 
      NEXT_REGISTERS_9_37_port, NEXT_REGISTERS_9_36_port, 
      NEXT_REGISTERS_9_35_port, NEXT_REGISTERS_9_34_port, 
      NEXT_REGISTERS_9_33_port, NEXT_REGISTERS_9_32_port, 
      NEXT_REGISTERS_9_31_port, NEXT_REGISTERS_9_30_port, 
      NEXT_REGISTERS_9_29_port, NEXT_REGISTERS_9_28_port, 
      NEXT_REGISTERS_9_27_port, NEXT_REGISTERS_9_26_port, 
      NEXT_REGISTERS_9_25_port, NEXT_REGISTERS_9_24_port, 
      NEXT_REGISTERS_9_23_port, NEXT_REGISTERS_9_22_port, 
      NEXT_REGISTERS_9_21_port, NEXT_REGISTERS_9_20_port, 
      NEXT_REGISTERS_9_19_port, NEXT_REGISTERS_9_18_port, 
      NEXT_REGISTERS_9_17_port, NEXT_REGISTERS_9_16_port, 
      NEXT_REGISTERS_9_15_port, NEXT_REGISTERS_9_14_port, 
      NEXT_REGISTERS_9_13_port, NEXT_REGISTERS_9_12_port, 
      NEXT_REGISTERS_9_11_port, NEXT_REGISTERS_9_10_port, 
      NEXT_REGISTERS_9_9_port, NEXT_REGISTERS_9_8_port, NEXT_REGISTERS_9_7_port
      , NEXT_REGISTERS_9_6_port, NEXT_REGISTERS_9_5_port, 
      NEXT_REGISTERS_9_4_port, NEXT_REGISTERS_9_3_port, NEXT_REGISTERS_9_2_port
      , NEXT_REGISTERS_9_1_port, NEXT_REGISTERS_9_0_port, 
      NEXT_REGISTERS_10_63_port, NEXT_REGISTERS_10_62_port, 
      NEXT_REGISTERS_10_61_port, NEXT_REGISTERS_10_60_port, 
      NEXT_REGISTERS_10_59_port, NEXT_REGISTERS_10_58_port, 
      NEXT_REGISTERS_10_57_port, NEXT_REGISTERS_10_56_port, 
      NEXT_REGISTERS_10_55_port, NEXT_REGISTERS_10_54_port, 
      NEXT_REGISTERS_10_53_port, NEXT_REGISTERS_10_52_port, 
      NEXT_REGISTERS_10_51_port, NEXT_REGISTERS_10_50_port, 
      NEXT_REGISTERS_10_49_port, NEXT_REGISTERS_10_48_port, 
      NEXT_REGISTERS_10_47_port, NEXT_REGISTERS_10_46_port, 
      NEXT_REGISTERS_10_45_port, NEXT_REGISTERS_10_44_port, 
      NEXT_REGISTERS_10_43_port, NEXT_REGISTERS_10_42_port, 
      NEXT_REGISTERS_10_41_port, NEXT_REGISTERS_10_40_port, 
      NEXT_REGISTERS_10_39_port, NEXT_REGISTERS_10_38_port, 
      NEXT_REGISTERS_10_37_port, NEXT_REGISTERS_10_36_port, 
      NEXT_REGISTERS_10_35_port, NEXT_REGISTERS_10_34_port, 
      NEXT_REGISTERS_10_33_port, NEXT_REGISTERS_10_32_port, 
      NEXT_REGISTERS_10_31_port, NEXT_REGISTERS_10_30_port, 
      NEXT_REGISTERS_10_29_port, NEXT_REGISTERS_10_28_port, 
      NEXT_REGISTERS_10_27_port, NEXT_REGISTERS_10_26_port, 
      NEXT_REGISTERS_10_25_port, NEXT_REGISTERS_10_24_port, 
      NEXT_REGISTERS_10_23_port, NEXT_REGISTERS_10_22_port, 
      NEXT_REGISTERS_10_21_port, NEXT_REGISTERS_10_20_port, 
      NEXT_REGISTERS_10_19_port, NEXT_REGISTERS_10_18_port, 
      NEXT_REGISTERS_10_17_port, NEXT_REGISTERS_10_16_port, 
      NEXT_REGISTERS_10_15_port, NEXT_REGISTERS_10_14_port, 
      NEXT_REGISTERS_10_13_port, NEXT_REGISTERS_10_12_port, 
      NEXT_REGISTERS_10_11_port, NEXT_REGISTERS_10_10_port, 
      NEXT_REGISTERS_10_9_port, NEXT_REGISTERS_10_8_port, 
      NEXT_REGISTERS_10_7_port, NEXT_REGISTERS_10_6_port, 
      NEXT_REGISTERS_10_5_port, NEXT_REGISTERS_10_4_port, 
      NEXT_REGISTERS_10_3_port, NEXT_REGISTERS_10_2_port, 
      NEXT_REGISTERS_10_1_port, NEXT_REGISTERS_10_0_port, 
      NEXT_REGISTERS_11_63_port, NEXT_REGISTERS_11_62_port, 
      NEXT_REGISTERS_11_61_port, NEXT_REGISTERS_11_60_port, 
      NEXT_REGISTERS_11_59_port, NEXT_REGISTERS_11_58_port, 
      NEXT_REGISTERS_11_57_port, NEXT_REGISTERS_11_56_port, 
      NEXT_REGISTERS_11_55_port, NEXT_REGISTERS_11_54_port, 
      NEXT_REGISTERS_11_53_port, NEXT_REGISTERS_11_52_port, 
      NEXT_REGISTERS_11_51_port, NEXT_REGISTERS_11_50_port, 
      NEXT_REGISTERS_11_49_port, NEXT_REGISTERS_11_48_port, 
      NEXT_REGISTERS_11_47_port, NEXT_REGISTERS_11_46_port, 
      NEXT_REGISTERS_11_45_port, NEXT_REGISTERS_11_44_port, 
      NEXT_REGISTERS_11_43_port, NEXT_REGISTERS_11_42_port, 
      NEXT_REGISTERS_11_41_port, NEXT_REGISTERS_11_40_port, 
      NEXT_REGISTERS_11_39_port, NEXT_REGISTERS_11_38_port, 
      NEXT_REGISTERS_11_37_port, NEXT_REGISTERS_11_36_port, 
      NEXT_REGISTERS_11_35_port, NEXT_REGISTERS_11_34_port, 
      NEXT_REGISTERS_11_33_port, NEXT_REGISTERS_11_32_port, 
      NEXT_REGISTERS_11_31_port, NEXT_REGISTERS_11_30_port, 
      NEXT_REGISTERS_11_29_port, NEXT_REGISTERS_11_28_port, 
      NEXT_REGISTERS_11_27_port, NEXT_REGISTERS_11_26_port, 
      NEXT_REGISTERS_11_25_port, NEXT_REGISTERS_11_24_port, 
      NEXT_REGISTERS_11_23_port, NEXT_REGISTERS_11_22_port, 
      NEXT_REGISTERS_11_21_port, NEXT_REGISTERS_11_20_port, 
      NEXT_REGISTERS_11_19_port, NEXT_REGISTERS_11_18_port, 
      NEXT_REGISTERS_11_17_port, NEXT_REGISTERS_11_16_port, 
      NEXT_REGISTERS_11_15_port, NEXT_REGISTERS_11_14_port, 
      NEXT_REGISTERS_11_13_port, NEXT_REGISTERS_11_12_port, 
      NEXT_REGISTERS_11_11_port, NEXT_REGISTERS_11_10_port, 
      NEXT_REGISTERS_11_9_port, NEXT_REGISTERS_11_8_port, 
      NEXT_REGISTERS_11_7_port, NEXT_REGISTERS_11_6_port, 
      NEXT_REGISTERS_11_5_port, NEXT_REGISTERS_11_4_port, 
      NEXT_REGISTERS_11_3_port, NEXT_REGISTERS_11_2_port, 
      NEXT_REGISTERS_11_1_port, NEXT_REGISTERS_11_0_port, 
      NEXT_REGISTERS_12_63_port, NEXT_REGISTERS_12_62_port, 
      NEXT_REGISTERS_12_61_port, NEXT_REGISTERS_12_60_port, 
      NEXT_REGISTERS_12_59_port, NEXT_REGISTERS_12_58_port, 
      NEXT_REGISTERS_12_57_port, NEXT_REGISTERS_12_56_port, 
      NEXT_REGISTERS_12_55_port, NEXT_REGISTERS_12_54_port, 
      NEXT_REGISTERS_12_53_port, NEXT_REGISTERS_12_52_port, 
      NEXT_REGISTERS_12_51_port, NEXT_REGISTERS_12_50_port, 
      NEXT_REGISTERS_12_49_port, NEXT_REGISTERS_12_48_port, 
      NEXT_REGISTERS_12_47_port, NEXT_REGISTERS_12_46_port, 
      NEXT_REGISTERS_12_45_port, NEXT_REGISTERS_12_44_port, 
      NEXT_REGISTERS_12_43_port, NEXT_REGISTERS_12_42_port, 
      NEXT_REGISTERS_12_41_port, NEXT_REGISTERS_12_40_port, 
      NEXT_REGISTERS_12_39_port, NEXT_REGISTERS_12_38_port, 
      NEXT_REGISTERS_12_37_port, NEXT_REGISTERS_12_36_port, 
      NEXT_REGISTERS_12_35_port, NEXT_REGISTERS_12_34_port, 
      NEXT_REGISTERS_12_33_port, NEXT_REGISTERS_12_32_port, 
      NEXT_REGISTERS_12_31_port, NEXT_REGISTERS_12_30_port, 
      NEXT_REGISTERS_12_29_port, NEXT_REGISTERS_12_28_port, 
      NEXT_REGISTERS_12_27_port, NEXT_REGISTERS_12_26_port, 
      NEXT_REGISTERS_12_25_port, NEXT_REGISTERS_12_24_port, 
      NEXT_REGISTERS_12_23_port, NEXT_REGISTERS_12_22_port, 
      NEXT_REGISTERS_12_21_port, NEXT_REGISTERS_12_20_port, 
      NEXT_REGISTERS_12_19_port, NEXT_REGISTERS_12_18_port, 
      NEXT_REGISTERS_12_17_port, NEXT_REGISTERS_12_16_port, 
      NEXT_REGISTERS_12_15_port, NEXT_REGISTERS_12_14_port, 
      NEXT_REGISTERS_12_13_port, NEXT_REGISTERS_12_12_port, 
      NEXT_REGISTERS_12_11_port, NEXT_REGISTERS_12_10_port, 
      NEXT_REGISTERS_12_9_port, NEXT_REGISTERS_12_8_port, 
      NEXT_REGISTERS_12_7_port, NEXT_REGISTERS_12_6_port, 
      NEXT_REGISTERS_12_5_port, NEXT_REGISTERS_12_4_port, 
      NEXT_REGISTERS_12_3_port, NEXT_REGISTERS_12_2_port, 
      NEXT_REGISTERS_12_1_port, NEXT_REGISTERS_12_0_port, 
      NEXT_REGISTERS_13_63_port, NEXT_REGISTERS_13_62_port, 
      NEXT_REGISTERS_13_61_port, NEXT_REGISTERS_13_60_port, 
      NEXT_REGISTERS_13_59_port, NEXT_REGISTERS_13_58_port, 
      NEXT_REGISTERS_13_57_port, NEXT_REGISTERS_13_56_port, 
      NEXT_REGISTERS_13_55_port, NEXT_REGISTERS_13_54_port, 
      NEXT_REGISTERS_13_53_port, NEXT_REGISTERS_13_52_port, 
      NEXT_REGISTERS_13_51_port, NEXT_REGISTERS_13_50_port, 
      NEXT_REGISTERS_13_49_port, NEXT_REGISTERS_13_48_port, 
      NEXT_REGISTERS_13_47_port, NEXT_REGISTERS_13_46_port, 
      NEXT_REGISTERS_13_45_port, NEXT_REGISTERS_13_44_port, 
      NEXT_REGISTERS_13_43_port, NEXT_REGISTERS_13_42_port, 
      NEXT_REGISTERS_13_41_port, NEXT_REGISTERS_13_40_port, 
      NEXT_REGISTERS_13_39_port, NEXT_REGISTERS_13_38_port, 
      NEXT_REGISTERS_13_37_port, NEXT_REGISTERS_13_36_port, 
      NEXT_REGISTERS_13_35_port, NEXT_REGISTERS_13_34_port, 
      NEXT_REGISTERS_13_33_port, NEXT_REGISTERS_13_32_port, 
      NEXT_REGISTERS_13_31_port, NEXT_REGISTERS_13_30_port, 
      NEXT_REGISTERS_13_29_port, NEXT_REGISTERS_13_28_port, 
      NEXT_REGISTERS_13_27_port, NEXT_REGISTERS_13_26_port, 
      NEXT_REGISTERS_13_25_port, NEXT_REGISTERS_13_24_port, 
      NEXT_REGISTERS_13_23_port, NEXT_REGISTERS_13_22_port, 
      NEXT_REGISTERS_13_21_port, NEXT_REGISTERS_13_20_port, 
      NEXT_REGISTERS_13_19_port, NEXT_REGISTERS_13_18_port, 
      NEXT_REGISTERS_13_17_port, NEXT_REGISTERS_13_16_port, 
      NEXT_REGISTERS_13_15_port, NEXT_REGISTERS_13_14_port, 
      NEXT_REGISTERS_13_13_port, NEXT_REGISTERS_13_12_port, 
      NEXT_REGISTERS_13_11_port, NEXT_REGISTERS_13_10_port, 
      NEXT_REGISTERS_13_9_port, NEXT_REGISTERS_13_8_port, 
      NEXT_REGISTERS_13_7_port, NEXT_REGISTERS_13_6_port, 
      NEXT_REGISTERS_13_5_port, NEXT_REGISTERS_13_4_port, 
      NEXT_REGISTERS_13_3_port, NEXT_REGISTERS_13_2_port, 
      NEXT_REGISTERS_13_1_port, NEXT_REGISTERS_13_0_port, 
      NEXT_REGISTERS_14_63_port, NEXT_REGISTERS_14_62_port, 
      NEXT_REGISTERS_14_61_port, NEXT_REGISTERS_14_60_port, 
      NEXT_REGISTERS_14_59_port, NEXT_REGISTERS_14_58_port, 
      NEXT_REGISTERS_14_57_port, NEXT_REGISTERS_14_56_port, 
      NEXT_REGISTERS_14_55_port, NEXT_REGISTERS_14_54_port, 
      NEXT_REGISTERS_14_53_port, NEXT_REGISTERS_14_52_port, 
      NEXT_REGISTERS_14_51_port, NEXT_REGISTERS_14_50_port, 
      NEXT_REGISTERS_14_49_port, NEXT_REGISTERS_14_48_port, 
      NEXT_REGISTERS_14_47_port, NEXT_REGISTERS_14_46_port, 
      NEXT_REGISTERS_14_45_port, NEXT_REGISTERS_14_44_port, 
      NEXT_REGISTERS_14_43_port, NEXT_REGISTERS_14_42_port, 
      NEXT_REGISTERS_14_41_port, NEXT_REGISTERS_14_40_port, 
      NEXT_REGISTERS_14_39_port, NEXT_REGISTERS_14_38_port, 
      NEXT_REGISTERS_14_37_port, NEXT_REGISTERS_14_36_port, 
      NEXT_REGISTERS_14_35_port, NEXT_REGISTERS_14_34_port, 
      NEXT_REGISTERS_14_33_port, NEXT_REGISTERS_14_32_port, 
      NEXT_REGISTERS_14_31_port, NEXT_REGISTERS_14_30_port, 
      NEXT_REGISTERS_14_29_port, NEXT_REGISTERS_14_28_port, 
      NEXT_REGISTERS_14_27_port, NEXT_REGISTERS_14_26_port, 
      NEXT_REGISTERS_14_25_port, NEXT_REGISTERS_14_24_port, 
      NEXT_REGISTERS_14_23_port, NEXT_REGISTERS_14_22_port, 
      NEXT_REGISTERS_14_21_port, NEXT_REGISTERS_14_20_port, 
      NEXT_REGISTERS_14_19_port, NEXT_REGISTERS_14_18_port, 
      NEXT_REGISTERS_14_17_port, NEXT_REGISTERS_14_16_port, 
      NEXT_REGISTERS_14_15_port, NEXT_REGISTERS_14_14_port, 
      NEXT_REGISTERS_14_13_port, NEXT_REGISTERS_14_12_port, 
      NEXT_REGISTERS_14_11_port, NEXT_REGISTERS_14_10_port, 
      NEXT_REGISTERS_14_9_port, NEXT_REGISTERS_14_8_port, 
      NEXT_REGISTERS_14_7_port, NEXT_REGISTERS_14_6_port, 
      NEXT_REGISTERS_14_5_port, NEXT_REGISTERS_14_4_port, 
      NEXT_REGISTERS_14_3_port, NEXT_REGISTERS_14_2_port, 
      NEXT_REGISTERS_14_1_port, NEXT_REGISTERS_14_0_port, 
      NEXT_REGISTERS_15_63_port, NEXT_REGISTERS_15_62_port, 
      NEXT_REGISTERS_15_61_port, NEXT_REGISTERS_15_60_port, 
      NEXT_REGISTERS_15_59_port, NEXT_REGISTERS_15_58_port, 
      NEXT_REGISTERS_15_57_port, NEXT_REGISTERS_15_56_port, 
      NEXT_REGISTERS_15_55_port, NEXT_REGISTERS_15_54_port, 
      NEXT_REGISTERS_15_53_port, NEXT_REGISTERS_15_52_port, 
      NEXT_REGISTERS_15_51_port, NEXT_REGISTERS_15_50_port, 
      NEXT_REGISTERS_15_49_port, NEXT_REGISTERS_15_48_port, 
      NEXT_REGISTERS_15_47_port, NEXT_REGISTERS_15_46_port, 
      NEXT_REGISTERS_15_45_port, NEXT_REGISTERS_15_44_port, 
      NEXT_REGISTERS_15_43_port, NEXT_REGISTERS_15_42_port, 
      NEXT_REGISTERS_15_41_port, NEXT_REGISTERS_15_40_port, 
      NEXT_REGISTERS_15_39_port, NEXT_REGISTERS_15_38_port, 
      NEXT_REGISTERS_15_37_port, NEXT_REGISTERS_15_36_port, 
      NEXT_REGISTERS_15_35_port, NEXT_REGISTERS_15_34_port, 
      NEXT_REGISTERS_15_33_port, NEXT_REGISTERS_15_32_port, 
      NEXT_REGISTERS_15_31_port, NEXT_REGISTERS_15_30_port, 
      NEXT_REGISTERS_15_29_port, NEXT_REGISTERS_15_28_port, 
      NEXT_REGISTERS_15_27_port, NEXT_REGISTERS_15_26_port, 
      NEXT_REGISTERS_15_25_port, NEXT_REGISTERS_15_24_port, 
      NEXT_REGISTERS_15_23_port, NEXT_REGISTERS_15_22_port, 
      NEXT_REGISTERS_15_21_port, NEXT_REGISTERS_15_20_port, 
      NEXT_REGISTERS_15_19_port, NEXT_REGISTERS_15_18_port, 
      NEXT_REGISTERS_15_17_port, NEXT_REGISTERS_15_16_port, 
      NEXT_REGISTERS_15_15_port, NEXT_REGISTERS_15_14_port, 
      NEXT_REGISTERS_15_13_port, NEXT_REGISTERS_15_12_port, 
      NEXT_REGISTERS_15_11_port, NEXT_REGISTERS_15_10_port, 
      NEXT_REGISTERS_15_9_port, NEXT_REGISTERS_15_8_port, 
      NEXT_REGISTERS_15_7_port, NEXT_REGISTERS_15_6_port, 
      NEXT_REGISTERS_15_5_port, NEXT_REGISTERS_15_4_port, 
      NEXT_REGISTERS_15_3_port, NEXT_REGISTERS_15_2_port, 
      NEXT_REGISTERS_15_1_port, NEXT_REGISTERS_15_0_port, 
      NEXT_REGISTERS_16_63_port, NEXT_REGISTERS_16_62_port, 
      NEXT_REGISTERS_16_61_port, NEXT_REGISTERS_16_60_port, 
      NEXT_REGISTERS_16_59_port, NEXT_REGISTERS_16_58_port, 
      NEXT_REGISTERS_16_57_port, NEXT_REGISTERS_16_56_port, 
      NEXT_REGISTERS_16_55_port, NEXT_REGISTERS_16_54_port, 
      NEXT_REGISTERS_16_53_port, NEXT_REGISTERS_16_52_port, 
      NEXT_REGISTERS_16_51_port, NEXT_REGISTERS_16_50_port, 
      NEXT_REGISTERS_16_49_port, NEXT_REGISTERS_16_48_port, 
      NEXT_REGISTERS_16_47_port, NEXT_REGISTERS_16_46_port, 
      NEXT_REGISTERS_16_45_port, NEXT_REGISTERS_16_44_port, 
      NEXT_REGISTERS_16_43_port, NEXT_REGISTERS_16_42_port, 
      NEXT_REGISTERS_16_41_port, NEXT_REGISTERS_16_40_port, 
      NEXT_REGISTERS_16_39_port, NEXT_REGISTERS_16_38_port, 
      NEXT_REGISTERS_16_37_port, NEXT_REGISTERS_16_36_port, 
      NEXT_REGISTERS_16_35_port, NEXT_REGISTERS_16_34_port, 
      NEXT_REGISTERS_16_33_port, NEXT_REGISTERS_16_32_port, 
      NEXT_REGISTERS_16_31_port, NEXT_REGISTERS_16_30_port, 
      NEXT_REGISTERS_16_29_port, NEXT_REGISTERS_16_28_port, 
      NEXT_REGISTERS_16_27_port, NEXT_REGISTERS_16_26_port, 
      NEXT_REGISTERS_16_25_port, NEXT_REGISTERS_16_24_port, 
      NEXT_REGISTERS_16_23_port, NEXT_REGISTERS_16_22_port, 
      NEXT_REGISTERS_16_21_port, NEXT_REGISTERS_16_20_port, 
      NEXT_REGISTERS_16_19_port, NEXT_REGISTERS_16_18_port, 
      NEXT_REGISTERS_16_17_port, NEXT_REGISTERS_16_16_port, 
      NEXT_REGISTERS_16_15_port, NEXT_REGISTERS_16_14_port, 
      NEXT_REGISTERS_16_13_port, NEXT_REGISTERS_16_12_port, 
      NEXT_REGISTERS_16_11_port, NEXT_REGISTERS_16_10_port, 
      NEXT_REGISTERS_16_9_port, NEXT_REGISTERS_16_8_port, 
      NEXT_REGISTERS_16_7_port, NEXT_REGISTERS_16_6_port, 
      NEXT_REGISTERS_16_5_port, NEXT_REGISTERS_16_4_port, 
      NEXT_REGISTERS_16_3_port, NEXT_REGISTERS_16_2_port, 
      NEXT_REGISTERS_16_1_port, NEXT_REGISTERS_16_0_port, 
      NEXT_REGISTERS_17_63_port, NEXT_REGISTERS_17_62_port, 
      NEXT_REGISTERS_17_61_port, NEXT_REGISTERS_17_60_port, 
      NEXT_REGISTERS_17_59_port, NEXT_REGISTERS_17_58_port, 
      NEXT_REGISTERS_17_57_port, NEXT_REGISTERS_17_56_port, 
      NEXT_REGISTERS_17_55_port, NEXT_REGISTERS_17_54_port, 
      NEXT_REGISTERS_17_53_port, NEXT_REGISTERS_17_52_port, 
      NEXT_REGISTERS_17_51_port, NEXT_REGISTERS_17_50_port, 
      NEXT_REGISTERS_17_49_port, NEXT_REGISTERS_17_48_port, 
      NEXT_REGISTERS_17_47_port, NEXT_REGISTERS_17_46_port, 
      NEXT_REGISTERS_17_45_port, NEXT_REGISTERS_17_44_port, 
      NEXT_REGISTERS_17_43_port, NEXT_REGISTERS_17_42_port, 
      NEXT_REGISTERS_17_41_port, NEXT_REGISTERS_17_40_port, 
      NEXT_REGISTERS_17_39_port, NEXT_REGISTERS_17_38_port, 
      NEXT_REGISTERS_17_37_port, NEXT_REGISTERS_17_36_port, 
      NEXT_REGISTERS_17_35_port, NEXT_REGISTERS_17_34_port, 
      NEXT_REGISTERS_17_33_port, NEXT_REGISTERS_17_32_port, 
      NEXT_REGISTERS_17_31_port, NEXT_REGISTERS_17_30_port, 
      NEXT_REGISTERS_17_29_port, NEXT_REGISTERS_17_28_port, 
      NEXT_REGISTERS_17_27_port, NEXT_REGISTERS_17_26_port, 
      NEXT_REGISTERS_17_25_port, NEXT_REGISTERS_17_24_port, 
      NEXT_REGISTERS_17_23_port, NEXT_REGISTERS_17_22_port, 
      NEXT_REGISTERS_17_21_port, NEXT_REGISTERS_17_20_port, 
      NEXT_REGISTERS_17_19_port, NEXT_REGISTERS_17_18_port, 
      NEXT_REGISTERS_17_17_port, NEXT_REGISTERS_17_16_port, 
      NEXT_REGISTERS_17_15_port, NEXT_REGISTERS_17_14_port, 
      NEXT_REGISTERS_17_13_port, NEXT_REGISTERS_17_12_port, 
      NEXT_REGISTERS_17_11_port, NEXT_REGISTERS_17_10_port, 
      NEXT_REGISTERS_17_9_port, NEXT_REGISTERS_17_8_port, 
      NEXT_REGISTERS_17_7_port, NEXT_REGISTERS_17_6_port, 
      NEXT_REGISTERS_17_5_port, NEXT_REGISTERS_17_4_port, 
      NEXT_REGISTERS_17_3_port, NEXT_REGISTERS_17_2_port, 
      NEXT_REGISTERS_17_1_port, NEXT_REGISTERS_17_0_port, 
      NEXT_REGISTERS_18_63_port, NEXT_REGISTERS_18_62_port, 
      NEXT_REGISTERS_18_61_port, NEXT_REGISTERS_18_60_port, 
      NEXT_REGISTERS_18_59_port, NEXT_REGISTERS_18_58_port, 
      NEXT_REGISTERS_18_57_port, NEXT_REGISTERS_18_56_port, 
      NEXT_REGISTERS_18_55_port, NEXT_REGISTERS_18_54_port, 
      NEXT_REGISTERS_18_53_port, NEXT_REGISTERS_18_52_port, 
      NEXT_REGISTERS_18_51_port, NEXT_REGISTERS_18_50_port, 
      NEXT_REGISTERS_18_49_port, NEXT_REGISTERS_18_48_port, 
      NEXT_REGISTERS_18_47_port, NEXT_REGISTERS_18_46_port, 
      NEXT_REGISTERS_18_45_port, NEXT_REGISTERS_18_44_port, 
      NEXT_REGISTERS_18_43_port, NEXT_REGISTERS_18_42_port, 
      NEXT_REGISTERS_18_41_port, NEXT_REGISTERS_18_40_port, 
      NEXT_REGISTERS_18_39_port, NEXT_REGISTERS_18_38_port, 
      NEXT_REGISTERS_18_37_port, NEXT_REGISTERS_18_36_port, 
      NEXT_REGISTERS_18_35_port, NEXT_REGISTERS_18_34_port, 
      NEXT_REGISTERS_18_33_port, NEXT_REGISTERS_18_32_port, 
      NEXT_REGISTERS_18_31_port, NEXT_REGISTERS_18_30_port, 
      NEXT_REGISTERS_18_29_port, NEXT_REGISTERS_18_28_port, 
      NEXT_REGISTERS_18_27_port, NEXT_REGISTERS_18_26_port, 
      NEXT_REGISTERS_18_25_port, NEXT_REGISTERS_18_24_port, 
      NEXT_REGISTERS_18_23_port, NEXT_REGISTERS_18_22_port, 
      NEXT_REGISTERS_18_21_port, NEXT_REGISTERS_18_20_port, 
      NEXT_REGISTERS_18_19_port, NEXT_REGISTERS_18_18_port, 
      NEXT_REGISTERS_18_17_port, NEXT_REGISTERS_18_16_port, 
      NEXT_REGISTERS_18_15_port, NEXT_REGISTERS_18_14_port, 
      NEXT_REGISTERS_18_13_port, NEXT_REGISTERS_18_12_port, 
      NEXT_REGISTERS_18_11_port, NEXT_REGISTERS_18_10_port, 
      NEXT_REGISTERS_18_9_port, NEXT_REGISTERS_18_8_port, 
      NEXT_REGISTERS_18_7_port, NEXT_REGISTERS_18_6_port, 
      NEXT_REGISTERS_18_5_port, NEXT_REGISTERS_18_4_port, 
      NEXT_REGISTERS_18_3_port, NEXT_REGISTERS_18_2_port, 
      NEXT_REGISTERS_18_1_port, NEXT_REGISTERS_18_0_port, 
      NEXT_REGISTERS_19_63_port, NEXT_REGISTERS_19_62_port, 
      NEXT_REGISTERS_19_61_port, NEXT_REGISTERS_19_60_port, 
      NEXT_REGISTERS_19_59_port, NEXT_REGISTERS_19_58_port, 
      NEXT_REGISTERS_19_57_port, NEXT_REGISTERS_19_56_port, 
      NEXT_REGISTERS_19_55_port, NEXT_REGISTERS_19_54_port, 
      NEXT_REGISTERS_19_53_port, NEXT_REGISTERS_19_52_port, 
      NEXT_REGISTERS_19_51_port, NEXT_REGISTERS_19_50_port, 
      NEXT_REGISTERS_19_49_port, NEXT_REGISTERS_19_48_port, 
      NEXT_REGISTERS_19_47_port, NEXT_REGISTERS_19_46_port, 
      NEXT_REGISTERS_19_45_port, NEXT_REGISTERS_19_44_port, 
      NEXT_REGISTERS_19_43_port, NEXT_REGISTERS_19_42_port, 
      NEXT_REGISTERS_19_41_port, NEXT_REGISTERS_19_40_port, 
      NEXT_REGISTERS_19_39_port, NEXT_REGISTERS_19_38_port, 
      NEXT_REGISTERS_19_37_port, NEXT_REGISTERS_19_36_port, 
      NEXT_REGISTERS_19_35_port, NEXT_REGISTERS_19_34_port, 
      NEXT_REGISTERS_19_33_port, NEXT_REGISTERS_19_32_port, 
      NEXT_REGISTERS_19_31_port, NEXT_REGISTERS_19_30_port, 
      NEXT_REGISTERS_19_29_port, NEXT_REGISTERS_19_28_port, 
      NEXT_REGISTERS_19_27_port, NEXT_REGISTERS_19_26_port, 
      NEXT_REGISTERS_19_25_port, NEXT_REGISTERS_19_24_port, 
      NEXT_REGISTERS_19_23_port, NEXT_REGISTERS_19_22_port, 
      NEXT_REGISTERS_19_21_port, NEXT_REGISTERS_19_20_port, 
      NEXT_REGISTERS_19_19_port, NEXT_REGISTERS_19_18_port, 
      NEXT_REGISTERS_19_17_port, NEXT_REGISTERS_19_16_port, 
      NEXT_REGISTERS_19_15_port, NEXT_REGISTERS_19_14_port, 
      NEXT_REGISTERS_19_13_port, NEXT_REGISTERS_19_12_port, 
      NEXT_REGISTERS_19_11_port, NEXT_REGISTERS_19_10_port, 
      NEXT_REGISTERS_19_9_port, NEXT_REGISTERS_19_8_port, 
      NEXT_REGISTERS_19_7_port, NEXT_REGISTERS_19_6_port, 
      NEXT_REGISTERS_19_5_port, NEXT_REGISTERS_19_4_port, 
      NEXT_REGISTERS_19_3_port, NEXT_REGISTERS_19_2_port, 
      NEXT_REGISTERS_19_1_port, NEXT_REGISTERS_19_0_port, 
      NEXT_REGISTERS_20_63_port, NEXT_REGISTERS_20_62_port, 
      NEXT_REGISTERS_20_61_port, NEXT_REGISTERS_20_60_port, 
      NEXT_REGISTERS_20_59_port, NEXT_REGISTERS_20_58_port, 
      NEXT_REGISTERS_20_57_port, NEXT_REGISTERS_20_56_port, 
      NEXT_REGISTERS_20_55_port, NEXT_REGISTERS_20_54_port, 
      NEXT_REGISTERS_20_53_port, NEXT_REGISTERS_20_52_port, 
      NEXT_REGISTERS_20_51_port, NEXT_REGISTERS_20_50_port, 
      NEXT_REGISTERS_20_49_port, NEXT_REGISTERS_20_48_port, 
      NEXT_REGISTERS_20_47_port, NEXT_REGISTERS_20_46_port, 
      NEXT_REGISTERS_20_45_port, NEXT_REGISTERS_20_44_port, 
      NEXT_REGISTERS_20_43_port, NEXT_REGISTERS_20_42_port, 
      NEXT_REGISTERS_20_41_port, NEXT_REGISTERS_20_40_port, 
      NEXT_REGISTERS_20_39_port, NEXT_REGISTERS_20_38_port, 
      NEXT_REGISTERS_20_37_port, NEXT_REGISTERS_20_36_port, 
      NEXT_REGISTERS_20_35_port, NEXT_REGISTERS_20_34_port, 
      NEXT_REGISTERS_20_33_port, NEXT_REGISTERS_20_32_port, 
      NEXT_REGISTERS_20_31_port, NEXT_REGISTERS_20_30_port, 
      NEXT_REGISTERS_20_29_port, NEXT_REGISTERS_20_28_port, 
      NEXT_REGISTERS_20_27_port, NEXT_REGISTERS_20_26_port, 
      NEXT_REGISTERS_20_25_port, NEXT_REGISTERS_20_24_port, 
      NEXT_REGISTERS_20_23_port, NEXT_REGISTERS_20_22_port, 
      NEXT_REGISTERS_20_21_port, NEXT_REGISTERS_20_20_port, 
      NEXT_REGISTERS_20_19_port, NEXT_REGISTERS_20_18_port, 
      NEXT_REGISTERS_20_17_port, NEXT_REGISTERS_20_16_port, 
      NEXT_REGISTERS_20_15_port, NEXT_REGISTERS_20_14_port, 
      NEXT_REGISTERS_20_13_port, NEXT_REGISTERS_20_12_port, 
      NEXT_REGISTERS_20_11_port, NEXT_REGISTERS_20_10_port, 
      NEXT_REGISTERS_20_9_port, NEXT_REGISTERS_20_8_port, 
      NEXT_REGISTERS_20_7_port, NEXT_REGISTERS_20_6_port, 
      NEXT_REGISTERS_20_5_port, NEXT_REGISTERS_20_4_port, 
      NEXT_REGISTERS_20_3_port, NEXT_REGISTERS_20_2_port, 
      NEXT_REGISTERS_20_1_port, NEXT_REGISTERS_20_0_port, 
      NEXT_REGISTERS_21_63_port, NEXT_REGISTERS_21_62_port, 
      NEXT_REGISTERS_21_61_port, NEXT_REGISTERS_21_60_port, 
      NEXT_REGISTERS_21_59_port, NEXT_REGISTERS_21_58_port, 
      NEXT_REGISTERS_21_57_port, NEXT_REGISTERS_21_56_port, 
      NEXT_REGISTERS_21_55_port, NEXT_REGISTERS_21_54_port, 
      NEXT_REGISTERS_21_53_port, NEXT_REGISTERS_21_52_port, 
      NEXT_REGISTERS_21_51_port, NEXT_REGISTERS_21_50_port, 
      NEXT_REGISTERS_21_49_port, NEXT_REGISTERS_21_48_port, 
      NEXT_REGISTERS_21_47_port, NEXT_REGISTERS_21_46_port, 
      NEXT_REGISTERS_21_45_port, NEXT_REGISTERS_21_44_port, 
      NEXT_REGISTERS_21_43_port, NEXT_REGISTERS_21_42_port, 
      NEXT_REGISTERS_21_41_port, NEXT_REGISTERS_21_40_port, 
      NEXT_REGISTERS_21_39_port, NEXT_REGISTERS_21_38_port, 
      NEXT_REGISTERS_21_37_port, NEXT_REGISTERS_21_36_port, 
      NEXT_REGISTERS_21_35_port, NEXT_REGISTERS_21_34_port, 
      NEXT_REGISTERS_21_33_port, NEXT_REGISTERS_21_32_port, 
      NEXT_REGISTERS_21_31_port, NEXT_REGISTERS_21_30_port, 
      NEXT_REGISTERS_21_29_port, NEXT_REGISTERS_21_28_port, 
      NEXT_REGISTERS_21_27_port, NEXT_REGISTERS_21_26_port, 
      NEXT_REGISTERS_21_25_port, NEXT_REGISTERS_21_24_port, 
      NEXT_REGISTERS_21_23_port, NEXT_REGISTERS_21_22_port, 
      NEXT_REGISTERS_21_21_port, NEXT_REGISTERS_21_20_port, 
      NEXT_REGISTERS_21_19_port, NEXT_REGISTERS_21_18_port, 
      NEXT_REGISTERS_21_17_port, NEXT_REGISTERS_21_16_port, 
      NEXT_REGISTERS_21_15_port, NEXT_REGISTERS_21_14_port, 
      NEXT_REGISTERS_21_13_port, NEXT_REGISTERS_21_12_port, 
      NEXT_REGISTERS_21_11_port, NEXT_REGISTERS_21_10_port, 
      NEXT_REGISTERS_21_9_port, NEXT_REGISTERS_21_8_port, 
      NEXT_REGISTERS_21_7_port, NEXT_REGISTERS_21_6_port, 
      NEXT_REGISTERS_21_5_port, NEXT_REGISTERS_21_4_port, 
      NEXT_REGISTERS_21_3_port, NEXT_REGISTERS_21_2_port, 
      NEXT_REGISTERS_21_1_port, NEXT_REGISTERS_21_0_port, 
      NEXT_REGISTERS_22_63_port, NEXT_REGISTERS_22_62_port, 
      NEXT_REGISTERS_22_61_port, NEXT_REGISTERS_22_60_port, 
      NEXT_REGISTERS_22_59_port, NEXT_REGISTERS_22_58_port, 
      NEXT_REGISTERS_22_57_port, NEXT_REGISTERS_22_56_port, 
      NEXT_REGISTERS_22_55_port, NEXT_REGISTERS_22_54_port, 
      NEXT_REGISTERS_22_53_port, NEXT_REGISTERS_22_52_port, 
      NEXT_REGISTERS_22_51_port, NEXT_REGISTERS_22_50_port, 
      NEXT_REGISTERS_22_49_port, NEXT_REGISTERS_22_48_port, 
      NEXT_REGISTERS_22_47_port, NEXT_REGISTERS_22_46_port, 
      NEXT_REGISTERS_22_45_port, NEXT_REGISTERS_22_44_port, 
      NEXT_REGISTERS_22_43_port, NEXT_REGISTERS_22_42_port, 
      NEXT_REGISTERS_22_41_port, NEXT_REGISTERS_22_40_port, 
      NEXT_REGISTERS_22_39_port, NEXT_REGISTERS_22_38_port, 
      NEXT_REGISTERS_22_37_port, NEXT_REGISTERS_22_36_port, 
      NEXT_REGISTERS_22_35_port, NEXT_REGISTERS_22_34_port, 
      NEXT_REGISTERS_22_33_port, NEXT_REGISTERS_22_32_port, 
      NEXT_REGISTERS_22_31_port, NEXT_REGISTERS_22_30_port, 
      NEXT_REGISTERS_22_29_port, NEXT_REGISTERS_22_28_port, 
      NEXT_REGISTERS_22_27_port, NEXT_REGISTERS_22_26_port, 
      NEXT_REGISTERS_22_25_port, NEXT_REGISTERS_22_24_port, 
      NEXT_REGISTERS_22_23_port, NEXT_REGISTERS_22_22_port, 
      NEXT_REGISTERS_22_21_port, NEXT_REGISTERS_22_20_port, 
      NEXT_REGISTERS_22_19_port, NEXT_REGISTERS_22_18_port, 
      NEXT_REGISTERS_22_17_port, NEXT_REGISTERS_22_16_port, 
      NEXT_REGISTERS_22_15_port, NEXT_REGISTERS_22_14_port, 
      NEXT_REGISTERS_22_13_port, NEXT_REGISTERS_22_12_port, 
      NEXT_REGISTERS_22_11_port, NEXT_REGISTERS_22_10_port, 
      NEXT_REGISTERS_22_9_port, NEXT_REGISTERS_22_8_port, 
      NEXT_REGISTERS_22_7_port, NEXT_REGISTERS_22_6_port, 
      NEXT_REGISTERS_22_5_port, NEXT_REGISTERS_22_4_port, 
      NEXT_REGISTERS_22_3_port, NEXT_REGISTERS_22_2_port, 
      NEXT_REGISTERS_22_1_port, NEXT_REGISTERS_22_0_port, 
      NEXT_REGISTERS_23_63_port, NEXT_REGISTERS_23_62_port, 
      NEXT_REGISTERS_23_61_port, NEXT_REGISTERS_23_60_port, 
      NEXT_REGISTERS_23_59_port, NEXT_REGISTERS_23_58_port, 
      NEXT_REGISTERS_23_57_port, NEXT_REGISTERS_23_56_port, 
      NEXT_REGISTERS_23_55_port, NEXT_REGISTERS_23_54_port, 
      NEXT_REGISTERS_23_53_port, NEXT_REGISTERS_23_52_port, 
      NEXT_REGISTERS_23_51_port, NEXT_REGISTERS_23_50_port, 
      NEXT_REGISTERS_23_49_port, NEXT_REGISTERS_23_48_port, 
      NEXT_REGISTERS_23_47_port, NEXT_REGISTERS_23_46_port, 
      NEXT_REGISTERS_23_45_port, NEXT_REGISTERS_23_44_port, 
      NEXT_REGISTERS_23_43_port, NEXT_REGISTERS_23_42_port, 
      NEXT_REGISTERS_23_41_port, NEXT_REGISTERS_23_40_port, 
      NEXT_REGISTERS_23_39_port, NEXT_REGISTERS_23_38_port, 
      NEXT_REGISTERS_23_37_port, NEXT_REGISTERS_23_36_port, 
      NEXT_REGISTERS_23_35_port, NEXT_REGISTERS_23_34_port, 
      NEXT_REGISTERS_23_33_port, NEXT_REGISTERS_23_32_port, 
      NEXT_REGISTERS_23_31_port, NEXT_REGISTERS_23_30_port, 
      NEXT_REGISTERS_23_29_port, NEXT_REGISTERS_23_28_port, 
      NEXT_REGISTERS_23_27_port, NEXT_REGISTERS_23_26_port, 
      NEXT_REGISTERS_23_25_port, NEXT_REGISTERS_23_24_port, 
      NEXT_REGISTERS_23_23_port, NEXT_REGISTERS_23_22_port, 
      NEXT_REGISTERS_23_21_port, NEXT_REGISTERS_23_20_port, 
      NEXT_REGISTERS_23_19_port, NEXT_REGISTERS_23_18_port, 
      NEXT_REGISTERS_23_17_port, NEXT_REGISTERS_23_16_port, 
      NEXT_REGISTERS_23_15_port, NEXT_REGISTERS_23_14_port, 
      NEXT_REGISTERS_23_13_port, NEXT_REGISTERS_23_12_port, 
      NEXT_REGISTERS_23_11_port, NEXT_REGISTERS_23_10_port, 
      NEXT_REGISTERS_23_9_port, NEXT_REGISTERS_23_8_port, 
      NEXT_REGISTERS_23_7_port, NEXT_REGISTERS_23_6_port, 
      NEXT_REGISTERS_23_5_port, NEXT_REGISTERS_23_4_port, 
      NEXT_REGISTERS_23_3_port, NEXT_REGISTERS_23_2_port, 
      NEXT_REGISTERS_23_1_port, NEXT_REGISTERS_23_0_port, 
      NEXT_REGISTERS_24_63_port, NEXT_REGISTERS_24_62_port, 
      NEXT_REGISTERS_24_61_port, NEXT_REGISTERS_24_60_port, 
      NEXT_REGISTERS_24_59_port, NEXT_REGISTERS_24_58_port, 
      NEXT_REGISTERS_24_57_port, NEXT_REGISTERS_24_56_port, 
      NEXT_REGISTERS_24_55_port, NEXT_REGISTERS_24_54_port, 
      NEXT_REGISTERS_24_53_port, NEXT_REGISTERS_24_52_port, 
      NEXT_REGISTERS_24_51_port, NEXT_REGISTERS_24_50_port, 
      NEXT_REGISTERS_24_49_port, NEXT_REGISTERS_24_48_port, 
      NEXT_REGISTERS_24_47_port, NEXT_REGISTERS_24_46_port, 
      NEXT_REGISTERS_24_45_port, NEXT_REGISTERS_24_44_port, 
      NEXT_REGISTERS_24_43_port, NEXT_REGISTERS_24_42_port, 
      NEXT_REGISTERS_24_41_port, NEXT_REGISTERS_24_40_port, 
      NEXT_REGISTERS_24_39_port, NEXT_REGISTERS_24_38_port, 
      NEXT_REGISTERS_24_37_port, NEXT_REGISTERS_24_36_port, 
      NEXT_REGISTERS_24_35_port, NEXT_REGISTERS_24_34_port, 
      NEXT_REGISTERS_24_33_port, NEXT_REGISTERS_24_32_port, 
      NEXT_REGISTERS_24_31_port, NEXT_REGISTERS_24_30_port, 
      NEXT_REGISTERS_24_29_port, NEXT_REGISTERS_24_28_port, 
      NEXT_REGISTERS_24_27_port, NEXT_REGISTERS_24_26_port, 
      NEXT_REGISTERS_24_25_port, NEXT_REGISTERS_24_24_port, 
      NEXT_REGISTERS_24_23_port, NEXT_REGISTERS_24_22_port, 
      NEXT_REGISTERS_24_21_port, NEXT_REGISTERS_24_20_port, 
      NEXT_REGISTERS_24_19_port, NEXT_REGISTERS_24_18_port, 
      NEXT_REGISTERS_24_17_port, NEXT_REGISTERS_24_16_port, 
      NEXT_REGISTERS_24_15_port, NEXT_REGISTERS_24_14_port, 
      NEXT_REGISTERS_24_13_port, NEXT_REGISTERS_24_12_port, 
      NEXT_REGISTERS_24_11_port, NEXT_REGISTERS_24_10_port, 
      NEXT_REGISTERS_24_9_port, NEXT_REGISTERS_24_8_port, 
      NEXT_REGISTERS_24_7_port, NEXT_REGISTERS_24_6_port, 
      NEXT_REGISTERS_24_5_port, NEXT_REGISTERS_24_4_port, 
      NEXT_REGISTERS_24_3_port, NEXT_REGISTERS_24_2_port, 
      NEXT_REGISTERS_24_1_port, NEXT_REGISTERS_24_0_port, 
      NEXT_REGISTERS_25_63_port, NEXT_REGISTERS_25_62_port, 
      NEXT_REGISTERS_25_61_port, NEXT_REGISTERS_25_60_port, 
      NEXT_REGISTERS_25_59_port, NEXT_REGISTERS_25_58_port, 
      NEXT_REGISTERS_25_57_port, NEXT_REGISTERS_25_56_port, 
      NEXT_REGISTERS_25_55_port, NEXT_REGISTERS_25_54_port, 
      NEXT_REGISTERS_25_53_port, NEXT_REGISTERS_25_52_port, 
      NEXT_REGISTERS_25_51_port, NEXT_REGISTERS_25_50_port, 
      NEXT_REGISTERS_25_49_port, NEXT_REGISTERS_25_48_port, 
      NEXT_REGISTERS_25_47_port, NEXT_REGISTERS_25_46_port, 
      NEXT_REGISTERS_25_45_port, NEXT_REGISTERS_25_44_port, 
      NEXT_REGISTERS_25_43_port, NEXT_REGISTERS_25_42_port, 
      NEXT_REGISTERS_25_41_port, NEXT_REGISTERS_25_40_port, 
      NEXT_REGISTERS_25_39_port, NEXT_REGISTERS_25_38_port, 
      NEXT_REGISTERS_25_37_port, NEXT_REGISTERS_25_36_port, 
      NEXT_REGISTERS_25_35_port, NEXT_REGISTERS_25_34_port, 
      NEXT_REGISTERS_25_33_port, NEXT_REGISTERS_25_32_port, 
      NEXT_REGISTERS_25_31_port, NEXT_REGISTERS_25_30_port, 
      NEXT_REGISTERS_25_29_port, NEXT_REGISTERS_25_28_port, 
      NEXT_REGISTERS_25_27_port, NEXT_REGISTERS_25_26_port, 
      NEXT_REGISTERS_25_25_port, NEXT_REGISTERS_25_24_port, 
      NEXT_REGISTERS_25_23_port, NEXT_REGISTERS_25_22_port, 
      NEXT_REGISTERS_25_21_port, NEXT_REGISTERS_25_20_port, 
      NEXT_REGISTERS_25_19_port, NEXT_REGISTERS_25_18_port, 
      NEXT_REGISTERS_25_17_port, NEXT_REGISTERS_25_16_port, 
      NEXT_REGISTERS_25_15_port, NEXT_REGISTERS_25_14_port, 
      NEXT_REGISTERS_25_13_port, NEXT_REGISTERS_25_12_port, 
      NEXT_REGISTERS_25_11_port, NEXT_REGISTERS_25_10_port, 
      NEXT_REGISTERS_25_9_port, NEXT_REGISTERS_25_8_port, 
      NEXT_REGISTERS_25_7_port, NEXT_REGISTERS_25_6_port, 
      NEXT_REGISTERS_25_5_port, NEXT_REGISTERS_25_4_port, 
      NEXT_REGISTERS_25_3_port, NEXT_REGISTERS_25_2_port, 
      NEXT_REGISTERS_25_1_port, NEXT_REGISTERS_25_0_port, 
      NEXT_REGISTERS_26_63_port, NEXT_REGISTERS_26_62_port, 
      NEXT_REGISTERS_26_61_port, NEXT_REGISTERS_26_60_port, 
      NEXT_REGISTERS_26_59_port, NEXT_REGISTERS_26_58_port, 
      NEXT_REGISTERS_26_57_port, NEXT_REGISTERS_26_56_port, 
      NEXT_REGISTERS_26_55_port, NEXT_REGISTERS_26_54_port, 
      NEXT_REGISTERS_26_53_port, NEXT_REGISTERS_26_52_port, 
      NEXT_REGISTERS_26_51_port, NEXT_REGISTERS_26_50_port, 
      NEXT_REGISTERS_26_49_port, NEXT_REGISTERS_26_48_port, 
      NEXT_REGISTERS_26_47_port, NEXT_REGISTERS_26_46_port, 
      NEXT_REGISTERS_26_45_port, NEXT_REGISTERS_26_44_port, 
      NEXT_REGISTERS_26_43_port, NEXT_REGISTERS_26_42_port, 
      NEXT_REGISTERS_26_41_port, NEXT_REGISTERS_26_40_port, 
      NEXT_REGISTERS_26_39_port, NEXT_REGISTERS_26_38_port, 
      NEXT_REGISTERS_26_37_port, NEXT_REGISTERS_26_36_port, 
      NEXT_REGISTERS_26_35_port, NEXT_REGISTERS_26_34_port, 
      NEXT_REGISTERS_26_33_port, NEXT_REGISTERS_26_32_port, 
      NEXT_REGISTERS_26_31_port, NEXT_REGISTERS_26_30_port, 
      NEXT_REGISTERS_26_29_port, NEXT_REGISTERS_26_28_port, 
      NEXT_REGISTERS_26_27_port, NEXT_REGISTERS_26_26_port, 
      NEXT_REGISTERS_26_25_port, NEXT_REGISTERS_26_24_port, 
      NEXT_REGISTERS_26_23_port, NEXT_REGISTERS_26_22_port, 
      NEXT_REGISTERS_26_21_port, NEXT_REGISTERS_26_20_port, 
      NEXT_REGISTERS_26_19_port, NEXT_REGISTERS_26_18_port, 
      NEXT_REGISTERS_26_17_port, NEXT_REGISTERS_26_16_port, 
      NEXT_REGISTERS_26_15_port, NEXT_REGISTERS_26_14_port, 
      NEXT_REGISTERS_26_13_port, NEXT_REGISTERS_26_12_port, 
      NEXT_REGISTERS_26_11_port, NEXT_REGISTERS_26_10_port, 
      NEXT_REGISTERS_26_9_port, NEXT_REGISTERS_26_8_port, 
      NEXT_REGISTERS_26_7_port, NEXT_REGISTERS_26_6_port, 
      NEXT_REGISTERS_26_5_port, NEXT_REGISTERS_26_4_port, 
      NEXT_REGISTERS_26_3_port, NEXT_REGISTERS_26_2_port, 
      NEXT_REGISTERS_26_1_port, NEXT_REGISTERS_26_0_port, 
      NEXT_REGISTERS_27_63_port, NEXT_REGISTERS_27_62_port, 
      NEXT_REGISTERS_27_61_port, NEXT_REGISTERS_27_60_port, 
      NEXT_REGISTERS_27_59_port, NEXT_REGISTERS_27_58_port, 
      NEXT_REGISTERS_27_57_port, NEXT_REGISTERS_27_56_port, 
      NEXT_REGISTERS_27_55_port, NEXT_REGISTERS_27_54_port, 
      NEXT_REGISTERS_27_53_port, NEXT_REGISTERS_27_52_port, 
      NEXT_REGISTERS_27_51_port, NEXT_REGISTERS_27_50_port, 
      NEXT_REGISTERS_27_49_port, NEXT_REGISTERS_27_48_port, 
      NEXT_REGISTERS_27_47_port, NEXT_REGISTERS_27_46_port, 
      NEXT_REGISTERS_27_45_port, NEXT_REGISTERS_27_44_port, 
      NEXT_REGISTERS_27_43_port, NEXT_REGISTERS_27_42_port, 
      NEXT_REGISTERS_27_41_port, NEXT_REGISTERS_27_40_port, 
      NEXT_REGISTERS_27_39_port, NEXT_REGISTERS_27_38_port, 
      NEXT_REGISTERS_27_37_port, NEXT_REGISTERS_27_36_port, 
      NEXT_REGISTERS_27_35_port, NEXT_REGISTERS_27_34_port, 
      NEXT_REGISTERS_27_33_port, NEXT_REGISTERS_27_32_port, 
      NEXT_REGISTERS_27_31_port, NEXT_REGISTERS_27_30_port, 
      NEXT_REGISTERS_27_29_port, NEXT_REGISTERS_27_28_port, 
      NEXT_REGISTERS_27_27_port, NEXT_REGISTERS_27_26_port, 
      NEXT_REGISTERS_27_25_port, NEXT_REGISTERS_27_24_port, 
      NEXT_REGISTERS_27_23_port, NEXT_REGISTERS_27_22_port, 
      NEXT_REGISTERS_27_21_port, NEXT_REGISTERS_27_20_port, 
      NEXT_REGISTERS_27_19_port, NEXT_REGISTERS_27_18_port, 
      NEXT_REGISTERS_27_17_port, NEXT_REGISTERS_27_16_port, 
      NEXT_REGISTERS_27_15_port, NEXT_REGISTERS_27_14_port, 
      NEXT_REGISTERS_27_13_port, NEXT_REGISTERS_27_12_port, 
      NEXT_REGISTERS_27_11_port, NEXT_REGISTERS_27_10_port, 
      NEXT_REGISTERS_27_9_port, NEXT_REGISTERS_27_8_port, 
      NEXT_REGISTERS_27_7_port, NEXT_REGISTERS_27_6_port, 
      NEXT_REGISTERS_27_5_port, NEXT_REGISTERS_27_4_port, 
      NEXT_REGISTERS_27_3_port, NEXT_REGISTERS_27_2_port, 
      NEXT_REGISTERS_27_1_port, NEXT_REGISTERS_27_0_port, 
      NEXT_REGISTERS_28_63_port, NEXT_REGISTERS_28_62_port, 
      NEXT_REGISTERS_28_61_port, NEXT_REGISTERS_28_60_port, 
      NEXT_REGISTERS_28_59_port, NEXT_REGISTERS_28_58_port, 
      NEXT_REGISTERS_28_57_port, NEXT_REGISTERS_28_56_port, 
      NEXT_REGISTERS_28_55_port, NEXT_REGISTERS_28_54_port, 
      NEXT_REGISTERS_28_53_port, NEXT_REGISTERS_28_52_port, 
      NEXT_REGISTERS_28_51_port, NEXT_REGISTERS_28_50_port, 
      NEXT_REGISTERS_28_49_port, NEXT_REGISTERS_28_48_port, 
      NEXT_REGISTERS_28_47_port, NEXT_REGISTERS_28_46_port, 
      NEXT_REGISTERS_28_45_port, NEXT_REGISTERS_28_44_port, 
      NEXT_REGISTERS_28_43_port, NEXT_REGISTERS_28_42_port, 
      NEXT_REGISTERS_28_41_port, NEXT_REGISTERS_28_40_port, 
      NEXT_REGISTERS_28_39_port, NEXT_REGISTERS_28_38_port, 
      NEXT_REGISTERS_28_37_port, NEXT_REGISTERS_28_36_port, 
      NEXT_REGISTERS_28_35_port, NEXT_REGISTERS_28_34_port, 
      NEXT_REGISTERS_28_33_port, NEXT_REGISTERS_28_32_port, 
      NEXT_REGISTERS_28_31_port, NEXT_REGISTERS_28_30_port, 
      NEXT_REGISTERS_28_29_port, NEXT_REGISTERS_28_28_port, 
      NEXT_REGISTERS_28_27_port, NEXT_REGISTERS_28_26_port, 
      NEXT_REGISTERS_28_25_port, NEXT_REGISTERS_28_24_port, 
      NEXT_REGISTERS_28_23_port, NEXT_REGISTERS_28_22_port, 
      NEXT_REGISTERS_28_21_port, NEXT_REGISTERS_28_20_port, 
      NEXT_REGISTERS_28_19_port, NEXT_REGISTERS_28_18_port, 
      NEXT_REGISTERS_28_17_port, NEXT_REGISTERS_28_16_port, 
      NEXT_REGISTERS_28_15_port, NEXT_REGISTERS_28_14_port, 
      NEXT_REGISTERS_28_13_port, NEXT_REGISTERS_28_12_port, 
      NEXT_REGISTERS_28_11_port, NEXT_REGISTERS_28_10_port, 
      NEXT_REGISTERS_28_9_port, NEXT_REGISTERS_28_8_port, 
      NEXT_REGISTERS_28_7_port, NEXT_REGISTERS_28_6_port, 
      NEXT_REGISTERS_28_5_port, NEXT_REGISTERS_28_4_port, 
      NEXT_REGISTERS_28_3_port, NEXT_REGISTERS_28_2_port, 
      NEXT_REGISTERS_28_1_port, NEXT_REGISTERS_28_0_port, 
      NEXT_REGISTERS_29_63_port, NEXT_REGISTERS_29_62_port, 
      NEXT_REGISTERS_29_61_port, NEXT_REGISTERS_29_60_port, 
      NEXT_REGISTERS_29_59_port, NEXT_REGISTERS_29_58_port, 
      NEXT_REGISTERS_29_57_port, NEXT_REGISTERS_29_56_port, 
      NEXT_REGISTERS_29_55_port, NEXT_REGISTERS_29_54_port, 
      NEXT_REGISTERS_29_53_port, NEXT_REGISTERS_29_52_port, 
      NEXT_REGISTERS_29_51_port, NEXT_REGISTERS_29_50_port, 
      NEXT_REGISTERS_29_49_port, NEXT_REGISTERS_29_48_port, 
      NEXT_REGISTERS_29_47_port, NEXT_REGISTERS_29_46_port, 
      NEXT_REGISTERS_29_45_port, NEXT_REGISTERS_29_44_port, 
      NEXT_REGISTERS_29_43_port, NEXT_REGISTERS_29_42_port, 
      NEXT_REGISTERS_29_41_port, NEXT_REGISTERS_29_40_port, 
      NEXT_REGISTERS_29_39_port, NEXT_REGISTERS_29_38_port, 
      NEXT_REGISTERS_29_37_port, NEXT_REGISTERS_29_36_port, 
      NEXT_REGISTERS_29_35_port, NEXT_REGISTERS_29_34_port, 
      NEXT_REGISTERS_29_33_port, NEXT_REGISTERS_29_32_port, 
      NEXT_REGISTERS_29_31_port, NEXT_REGISTERS_29_30_port, 
      NEXT_REGISTERS_29_29_port, NEXT_REGISTERS_29_28_port, 
      NEXT_REGISTERS_29_27_port, NEXT_REGISTERS_29_26_port, 
      NEXT_REGISTERS_29_25_port, NEXT_REGISTERS_29_24_port, 
      NEXT_REGISTERS_29_23_port, NEXT_REGISTERS_29_22_port, 
      NEXT_REGISTERS_29_21_port, NEXT_REGISTERS_29_20_port, 
      NEXT_REGISTERS_29_19_port, NEXT_REGISTERS_29_18_port, 
      NEXT_REGISTERS_29_17_port, NEXT_REGISTERS_29_16_port, 
      NEXT_REGISTERS_29_15_port, NEXT_REGISTERS_29_14_port, 
      NEXT_REGISTERS_29_13_port, NEXT_REGISTERS_29_12_port, 
      NEXT_REGISTERS_29_11_port, NEXT_REGISTERS_29_10_port, 
      NEXT_REGISTERS_29_9_port, NEXT_REGISTERS_29_8_port, 
      NEXT_REGISTERS_29_7_port, NEXT_REGISTERS_29_6_port, 
      NEXT_REGISTERS_29_5_port, NEXT_REGISTERS_29_4_port, 
      NEXT_REGISTERS_29_3_port, NEXT_REGISTERS_29_2_port, 
      NEXT_REGISTERS_29_1_port, NEXT_REGISTERS_29_0_port, 
      NEXT_REGISTERS_30_63_port, NEXT_REGISTERS_30_62_port, 
      NEXT_REGISTERS_30_61_port, NEXT_REGISTERS_30_60_port, 
      NEXT_REGISTERS_30_59_port, NEXT_REGISTERS_30_58_port, 
      NEXT_REGISTERS_30_57_port, NEXT_REGISTERS_30_56_port, 
      NEXT_REGISTERS_30_55_port, NEXT_REGISTERS_30_54_port, 
      NEXT_REGISTERS_30_53_port, NEXT_REGISTERS_30_52_port, 
      NEXT_REGISTERS_30_51_port, NEXT_REGISTERS_30_50_port, 
      NEXT_REGISTERS_30_49_port, NEXT_REGISTERS_30_48_port, 
      NEXT_REGISTERS_30_47_port, NEXT_REGISTERS_30_46_port, 
      NEXT_REGISTERS_30_45_port, NEXT_REGISTERS_30_44_port, 
      NEXT_REGISTERS_30_43_port, NEXT_REGISTERS_30_42_port, 
      NEXT_REGISTERS_30_41_port, NEXT_REGISTERS_30_40_port, 
      NEXT_REGISTERS_30_39_port, NEXT_REGISTERS_30_38_port, 
      NEXT_REGISTERS_30_37_port, NEXT_REGISTERS_30_36_port, 
      NEXT_REGISTERS_30_35_port, NEXT_REGISTERS_30_34_port, 
      NEXT_REGISTERS_30_33_port, NEXT_REGISTERS_30_32_port, 
      NEXT_REGISTERS_30_31_port, NEXT_REGISTERS_30_30_port, 
      NEXT_REGISTERS_30_29_port, NEXT_REGISTERS_30_28_port, 
      NEXT_REGISTERS_30_27_port, NEXT_REGISTERS_30_26_port, 
      NEXT_REGISTERS_30_25_port, NEXT_REGISTERS_30_24_port, 
      NEXT_REGISTERS_30_23_port, NEXT_REGISTERS_30_22_port, 
      NEXT_REGISTERS_30_21_port, NEXT_REGISTERS_30_20_port, 
      NEXT_REGISTERS_30_19_port, NEXT_REGISTERS_30_18_port, 
      NEXT_REGISTERS_30_17_port, NEXT_REGISTERS_30_16_port, 
      NEXT_REGISTERS_30_15_port, NEXT_REGISTERS_30_14_port, 
      NEXT_REGISTERS_30_13_port, NEXT_REGISTERS_30_12_port, 
      NEXT_REGISTERS_30_11_port, NEXT_REGISTERS_30_10_port, 
      NEXT_REGISTERS_30_9_port, NEXT_REGISTERS_30_8_port, 
      NEXT_REGISTERS_30_7_port, NEXT_REGISTERS_30_6_port, 
      NEXT_REGISTERS_30_5_port, NEXT_REGISTERS_30_4_port, 
      NEXT_REGISTERS_30_3_port, NEXT_REGISTERS_30_2_port, 
      NEXT_REGISTERS_30_1_port, NEXT_REGISTERS_30_0_port, 
      NEXT_REGISTERS_31_63_port, NEXT_REGISTERS_31_62_port, 
      NEXT_REGISTERS_31_61_port, NEXT_REGISTERS_31_60_port, 
      NEXT_REGISTERS_31_59_port, NEXT_REGISTERS_31_58_port, 
      NEXT_REGISTERS_31_57_port, NEXT_REGISTERS_31_56_port, 
      NEXT_REGISTERS_31_55_port, NEXT_REGISTERS_31_54_port, 
      NEXT_REGISTERS_31_53_port, NEXT_REGISTERS_31_52_port, 
      NEXT_REGISTERS_31_51_port, NEXT_REGISTERS_31_50_port, 
      NEXT_REGISTERS_31_49_port, NEXT_REGISTERS_31_48_port, 
      NEXT_REGISTERS_31_47_port, NEXT_REGISTERS_31_46_port, 
      NEXT_REGISTERS_31_45_port, NEXT_REGISTERS_31_44_port, 
      NEXT_REGISTERS_31_43_port, NEXT_REGISTERS_31_42_port, 
      NEXT_REGISTERS_31_41_port, NEXT_REGISTERS_31_40_port, 
      NEXT_REGISTERS_31_39_port, NEXT_REGISTERS_31_38_port, 
      NEXT_REGISTERS_31_37_port, NEXT_REGISTERS_31_36_port, 
      NEXT_REGISTERS_31_35_port, NEXT_REGISTERS_31_34_port, 
      NEXT_REGISTERS_31_33_port, NEXT_REGISTERS_31_32_port, 
      NEXT_REGISTERS_31_31_port, NEXT_REGISTERS_31_30_port, 
      NEXT_REGISTERS_31_29_port, NEXT_REGISTERS_31_28_port, 
      NEXT_REGISTERS_31_27_port, NEXT_REGISTERS_31_26_port, 
      NEXT_REGISTERS_31_25_port, NEXT_REGISTERS_31_24_port, 
      NEXT_REGISTERS_31_23_port, NEXT_REGISTERS_31_22_port, 
      NEXT_REGISTERS_31_21_port, NEXT_REGISTERS_31_20_port, 
      NEXT_REGISTERS_31_19_port, NEXT_REGISTERS_31_18_port, 
      NEXT_REGISTERS_31_17_port, NEXT_REGISTERS_31_16_port, 
      NEXT_REGISTERS_31_15_port, NEXT_REGISTERS_31_14_port, 
      NEXT_REGISTERS_31_13_port, NEXT_REGISTERS_31_12_port, 
      NEXT_REGISTERS_31_11_port, NEXT_REGISTERS_31_10_port, 
      NEXT_REGISTERS_31_9_port, NEXT_REGISTERS_31_8_port, 
      NEXT_REGISTERS_31_7_port, NEXT_REGISTERS_31_6_port, 
      NEXT_REGISTERS_31_5_port, NEXT_REGISTERS_31_4_port, 
      NEXT_REGISTERS_31_3_port, NEXT_REGISTERS_31_2_port, 
      NEXT_REGISTERS_31_1_port, NEXT_REGISTERS_31_0_port, N22, N23, N24, N25, 
      N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40
      , N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, 
      N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69
      , N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, 
      N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98
      , N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, 
      N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, 
      N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, 
      N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
      N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
      N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, 
      N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, 
      N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, 
      N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, 
      N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, 
      N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, 
      N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, 
      N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, 
      N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, 
      N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, 
      N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, 
      N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, 
      N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, 
      N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, 
      N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, 
      N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, 
      N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, 
      N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, 
      N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, 
      N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, 
      N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, 
      N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, 
      N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, 
      N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, 
      N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, 
      N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, 
      N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, 
      N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, 
      N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, 
      N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, 
      N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, 
      N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, 
      N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, 
      N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, 
      N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, 
      N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, 
      N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, 
      N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, 
      N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, 
      N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, 
      N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, 
      N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, 
      N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, 
      N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, 
      N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, 
      N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, 
      N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, 
      N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, 
      N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, 
      N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, 
      N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, 
      N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, 
      N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, 
      N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, 
      N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, 
      N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, 
      N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, 
      N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, 
      N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, 
      N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, 
      N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, 
      N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, 
      N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, 
      N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, 
      N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, 
      N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, 
      N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, 
      N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, 
      N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, 
      N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, 
      N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, 
      N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, 
      N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, 
      N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, 
      N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, 
      N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, 
      N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, 
      N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, 
      N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, 
      N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, 
      N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, 
      N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, 
      N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, 
      N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, 
      N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, 
      N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, 
      N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, 
      N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, 
      N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, 
      N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, 
      N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, 
      N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, 
      N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, 
      N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, 
      N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, 
      N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, 
      N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, 
      N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, 
      N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, 
      N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, 
      N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, 
      N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, 
      N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, 
      N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, 
      N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, 
      N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, 
      N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, 
      N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, 
      N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, 
      N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, 
      N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, 
      N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, 
      N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, 
      N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, 
      N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, 
      N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, 
      N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, 
      N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, 
      N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, 
      N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, 
      N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, 
      N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, 
      N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, 
      N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, 
      N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, 
      N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, 
      N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, 
      N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, 
      N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, 
      N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, 
      N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, 
      N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, 
      N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, 
      N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, 
      N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, 
      N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, 
      N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, 
      N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, 
      N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, 
      N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, 
      N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718, 
      N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, 
      N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, 
      N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, 
      N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, 
      N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, 
      N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, 
      N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, 
      N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, 
      N1799, N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, 
      N1809, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, 
      N1819, N1820, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, 
      N1829, N1830, N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, 
      N1839, N1840, N1841, N1842, N1843, N1844, N1845, N1846, N1847, N1848, 
      N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, 
      N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, 
      N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, 
      N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1886, N1887, N1888, 
      N1889, N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, 
      N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, 
      N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, 
      N1919, N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, 
      N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, 
      N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, 
      N1949, N1950, N1951, N1952, N1953, N1954, N1955, N1956, N1957, N1958, 
      N1959, N1960, N1961, N1962, N1963, N1964, N1965, N1966, N1967, N1968, 
      N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1978, 
      N1979, N1980, N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1988, 
      N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, 
      N1999, N2000, N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, 
      N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, 
      N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, 
      N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, 
      N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, 
      N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, 
      N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, 
      N2069, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, 
      N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, 
      N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, 
      N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, 
      N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119, 
      N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2129, 
      N2130, N2131, N2132, N2133, N2134, N2136, N2137, N2138, N2139, N2140, 
      N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, 
      N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2159, N2160, 
      N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168, N2169, N2170, 
      N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2179, N2180, 
      N2181, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189, N2190, 
      N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199, N2234, 
      N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, 
      N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, 
      N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, 
      N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274, 
      N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, 
      N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294, 
      N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, 
      N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, 
      N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, 
      N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, 
      N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, 
      N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, 
      N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, 
      N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, 
      N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, 
      N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, 
      N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, 
      N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, 
      N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, 
      N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, 
      N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, 
      N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454, 
      N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464, 
      N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474, 
      N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, 
      N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, 
      N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, 
      N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, 
      N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, 
      N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, 
      N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, 
      N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, 
      N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564, 
      N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574, 
      N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584, 
      N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594, 
      N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, 
      N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, 
      N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, 
      N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, 
      N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, 
      N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, 
      N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, 
      N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, 
      N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, 
      N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, 
      N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, 
      N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714, 
      N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724, 
      N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734, 
      N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, 
      N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, 
      N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, 
      N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, 
      N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, 
      N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, 
      N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, 
      N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, 
      N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, 
      N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, 
      N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, 
      N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, 
      N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, 
      N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, 
      N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, 
      N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, 
      N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, 
      N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, 
      N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, 
      N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, 
      N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, 
      N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, 
      N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, 
      N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, 
      N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, 
      N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, 
      N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, 
      N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, 
      N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, 
      N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, 
      N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, 
      N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, 
      N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, 
      N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, 
      N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, 
      N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, 
      N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, 
      N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, 
      N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, 
      N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, 
      N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, 
      N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, 
      N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, 
      N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, 
      N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, 
      N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, 
      N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, 
      N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, 
      N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, 
      N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, 
      N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, 
      N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, 
      N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, 
      N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, 
      N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, 
      N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, 
      N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, 
      N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, 
      N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, 
      N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, 
      N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, 
      N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, 
      N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, 
      N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, 
      N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, 
      N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, 
      N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, 
      N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, 
      N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424, 
      N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434, 
      N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N3444, 
      N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, 
      N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464, 
      N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3474, 
      N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484, 
      N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, 
      N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, 
      N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, 
      N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, 
      N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, 
      N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, 
      N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554, 
      N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564, 
      N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574, 
      N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584, 
      N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594, 
      N3595, N3596, N3597, N3598, N3599, N3600, N3601, N3602, N3603, N3604, 
      N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614, 
      N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, 
      N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, 
      N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, 
      N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, 
      N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, 
      N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, 
      N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, 
      N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, 
      N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, 
      N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714, 
      N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, 
      N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, 
      N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744, 
      N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, 
      N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, 
      N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774, 
      N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, 
      N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, 
      N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, 
      N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, 
      N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824, 
      N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834, 
      N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3843, N3844, 
      N3845, N3846, N3847, N3848, N3849, N3850, N3851, N3852, N3853, N3854, 
      N3855, N3856, N3857, N3858, N3859, N3860, N3861, N3862, N3863, N3864, 
      N3865, N3866, N3867, N3868, N3869, N3870, N3871, N3872, N3873, N3874, 
      N3875, N3876, N3877, N3878, N3879, N3880, N3881, N3882, N3883, N3884, 
      N3885, N3886, N3887, N3888, N3889, N3890, N3891, N3892, N3893, N3894, 
      N3895, N3896, N3897, N3898, N3899, N3900, N3901, N3902, N3903, N3904, 
      N3905, N3906, N3907, N3908, N3909, N3910, N3911, N3912, N3913, N3914, 
      N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3922, N3923, N3924, 
      N3925, N3926, N3927, N3928, N3929, N3930, N3931, N3932, N3933, N3934, 
      N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944, 
      N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, 
      N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, 
      N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, 
      N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, 
      N3985, N3986, N3987, N3988, N3989, N3990, N3991, N3992, N3993, N3994, 
      N3995, N3996, N3997, N3998, N3999, N4000, N4001, N4002, N4003, N4004, 
      N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, 
      N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4022, N4023, N4024, 
      N4025, N4026, N4027, N4028, N4029, N4030, N4031, N4032, N4033, N4034, 
      N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4043, N4044, 
      N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054, 
      N4055, N4056, N4057, N4058, N4059, N4060, N4061, N4062, N4063, N4064, 
      N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073, N4074, 
      N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083, N4084, 
      N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093, N4094, 
      N4095, N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104, 
      N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114, 
      N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124, 
      N4125, N4126, N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134, 
      N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144, 
      N4145, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154, 
      N4155, N4156, N4157, N4158, N4159, N4160, N4161, N4162, N4163, N4164, 
      N4165, N4166, N4167, N4168, N4169, N4170, N4171, N4172, N4173, N4174, 
      N4175, N4176, N4177, N4178, N4179, N4180, N4181, N4182, N4183, N4184, 
      N4185, N4186, N4187, N4188, N4189, N4190, N4191, N4192, N4193, N4194, 
      N4195, N4196, N4197, N4198, N4199, N4200, N4201, N4202, N4203, N4204, 
      N4205, N4206, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214, 
      N4215, N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, 
      N4225, N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, 
      N4235, N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, 
      N4245, N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254, 
      N4255, N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264, 
      N4265, N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274, 
      N4275, N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, 
      N4285, N4286, N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294, 
      N4295, N4296, N4297, N4298, N4299, N4300, N4301, N4302, N4303, N4304, 
      N4305, N4306, N4307, N4308, N4309, N4310, N4311, N4312, N4313, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22_port, n23_port, n24_port, n25_port, n26_port, n27_port
      , n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, n34_port, 
      n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, n41_port, 
      n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, 
      n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, 
      n70_port, n71_port, n72_port, n73_port, n74_port, n75_port, n76_port, 
      n77_port, n78_port, n79_port, n80_port, n81_port, n82_port, n83_port, 
      n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, 
      n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, 
      n98_port, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port
      , n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114_port, n115_port, n116_port, 
      n117_port, n118_port, n119_port, n120_port, n121_port, n122_port, 
      n123_port, n124_port, n125_port, n126_port, n127_port, n128_port, 
      n129_port, n130_port, n131_port, n132_port, n133_port, n134_port, 
      n135_port, n136_port, n137_port, n138_port, n139_port, n140_port, 
      n141_port, n142_port, n143_port, n144_port, n145_port, n146_port, 
      n147_port, n148_port, n149_port, n150_port, n151_port, n152_port, 
      n153_port, n154_port, n155_port, n156_port, n157_port, n158_port, 
      n159_port, n160_port, n161_port, n162_port, n163_port, n164_port, 
      n165_port, n166_port, n167_port, n168_port, n169_port, n170_port, 
      n171_port, n172_port, n173_port, n174_port, n175_port, n176_port, 
      n177_port, n178_port, n179_port, n180_port, n181_port, n182_port, 
      n183_port, n184_port, n185_port, n186_port, n187_port, n188_port, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204_port, n205_port, n206_port, 
      n207_port, n208_port, n209_port, n210_port, n211_port, n212_port, 
      n213_port, n214_port, n215_port, n216_port, n217_port, n218_port, 
      n219_port, n220_port, n221_port, n222_port, n223_port, n224_port, 
      n225_port, n226_port, n227_port, n228_port, n229_port, n230_port, 
      n231_port, n232_port, n233_port, n234_port, n235_port, n236_port, 
      n237_port, n238_port, n239_port, n240_port, n241_port, n242_port, 
      n243_port, n244_port, n245_port, n246_port, n247_port, n248_port, 
      n249_port, n250_port, n251_port, n252_port, n253_port, n254_port, 
      n255_port, n256_port, n257_port, n258_port, n259_port, n260_port, 
      n261_port, n262_port, n263_port, n264_port, n265_port, n266_port, 
      n267_port, n268_port, n269_port, n270_port, n271_port, n272_port, 
      n273_port, n274_port, n275_port, n276_port, n277_port, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, 
      n285_port, n286_port, n287_port, n288_port, n289_port, n290_port, 
      n291_port, n292_port, n293_port, n294_port, n295_port, n296_port, 
      n297_port, n298_port, n299_port, n300_port, n301_port, n302_port, 
      n303_port, n304_port, n305_port, n306_port, n307_port, n308_port, 
      n309_port, n310_port, n311_port, n312_port, n313_port, n314_port, 
      n315_port, n316_port, n317_port, n318_port, n319_port, n320_port, 
      n321_port, n322_port, n323_port, n324_port, n325_port, n326_port, 
      n327_port, n328_port, n329_port, n330_port, n331_port, n332_port, 
      n333_port, n334_port, n335_port, n336_port, n337_port, n338_port, 
      n339_port, n340_port, n341_port, n342_port, n343_port, n344_port, 
      n345_port, n346_port, n347_port, n348_port, n349_port, n350_port, 
      n351_port, n352_port, n353_port, n354_port, n355_port, n356_port, 
      n357_port, n358_port, n359_port, n360_port, n361_port, n362_port, 
      n363_port, n364_port, n365_port, n366_port, n367_port, n368_port, 
      n369_port, n370_port, n371_port, n372_port, n373_port, n374_port, 
      n375_port, n376_port, n377_port, n378_port, n379_port, n380_port, 
      n381_port, n382_port, n383_port, n384_port, n385_port, n386_port, 
      n387_port, n388_port, n389_port, n390_port, n391_port, n392_port, 
      n393_port, n394_port, n395_port, n396_port, n397_port, n398_port, 
      n399_port, n400_port, n401_port, n402_port, n403_port, n404_port, 
      n405_port, n406_port, n407_port, n408_port, n409_port, n410_port, 
      n411_port, n412_port, n413_port, n414_port, n415_port, n416_port, 
      n417_port, n418_port, n419_port, n420_port, n421_port, n422_port, 
      n423_port, n424_port, n425_port, n426_port, n427_port, n428_port, 
      n429_port, n430_port, n431_port, n432_port, n433_port, n434_port, 
      n435_port, n436_port, n437_port, n438_port, n439_port, n440_port, 
      n441_port, n442_port, n443_port, n444_port, n445_port, n446_port, 
      n447_port, n448_port, n449_port, n450_port, n451_port, n452_port, 
      n453_port, n454_port, n455_port, n456_port, n457_port, n458_port, 
      n459_port, n460_port, n461_port, n462_port, n463_port, n464_port, 
      n465_port, n466_port, n467_port, n468_port, n469_port, n470_port, 
      n471_port, n472_port, n473_port, n474_port, n475_port, n476_port, 
      n477_port, n478_port, n479_port, n480_port, n481_port, n482_port, 
      n483_port, n484_port, n485_port, n486_port, n487_port, n488_port, 
      n489_port, n490_port, n491_port, n492_port, n493_port, n494_port, 
      n495_port, n496_port, n497_port, n498_port, n499_port, n500_port, 
      n501_port, n502_port, n503_port, n504_port, n505_port, n506_port, 
      n507_port, n508_port, n509_port, n510_port, n511_port, n512_port, 
      n513_port, n514_port, n515_port, n516_port, n517_port, n518_port, 
      n519_port, n520_port, n521_port, n522_port, n523_port, n524_port, 
      n525_port, n526_port, n527_port, n528_port, n529_port, n530_port, 
      n531_port, n532_port, n533_port, n534_port, n535_port, n536_port, 
      n537_port, n538_port, n539_port, n540_port, n541_port, n542_port, 
      n543_port, n544_port, n545_port, n546_port, n547_port, n548_port, 
      n549_port, n550_port, n551_port, n552_port, n553_port, n554_port, 
      n555_port, n556_port, n557_port, n558_port, n559_port, n560_port, 
      n561_port, n562_port, n563_port, n564_port, n565_port, n566_port, 
      n567_port, n568_port, n569_port, n570_port, n571_port, n572_port, 
      n573_port, n574_port, n575_port, n576_port, n577_port, n578_port, 
      n579_port, n580_port, n581_port, n582_port, n583_port, n584_port, 
      n585_port, n586_port, n587_port, n588_port, n589_port, n590_port, 
      n591_port, n592_port, n593_port, n594_port, n595_port, n596_port, 
      n597_port, n598_port, n599_port, n600_port, n601_port, n602_port, 
      n603_port, n604_port, n605_port, n606_port, n607_port, n608_port, 
      n609_port, n610_port, n611_port, n612_port, n613_port, n614_port, 
      n615_port, n616_port, n617_port, n618_port, n619_port, n620_port, 
      n621_port, n622_port, n623_port, n624_port, n625_port, n626_port, 
      n627_port, n628_port, n629_port, n630_port, n631_port, n632_port, 
      n633_port, n634_port, n635_port, n636_port, n637_port, n638_port, 
      n639_port, n640_port, n641_port, n642_port, n643_port, n644_port, 
      n645_port, n646_port, n647_port, n648_port, n649_port, n650_port, 
      n651_port, n652_port, n653_port, n654_port, n655_port, n656_port, 
      n657_port, n658_port, n659_port, n660_port, n661_port, n662_port, 
      n663_port, n664_port, n665_port, n666_port, n667_port, n668_port, 
      n669_port, n670_port, n671_port, n672_port, n673_port, n674_port, 
      n675_port, n676_port, n677_port, n678_port, n679_port, n680_port, 
      n681_port, n682_port, n683_port, n684_port, n685_port, n686_port, 
      n687_port, n688_port, n689_port, n690_port, n691_port, n692_port, 
      n693_port, n694_port, n695_port, n696_port, n697_port, n698_port, 
      n699_port, n700_port, n701_port, n702_port, n703_port, n704_port, 
      n705_port, n706_port, n707_port, n708_port, n709_port, n710_port, 
      n711_port, n712_port, n713_port, n714_port, n715_port, n716_port, 
      n717_port, n718_port, n719_port, n720_port, n721_port, n722_port, 
      n723_port, n724_port, n725_port, n726_port, n727_port, n728_port, 
      n729_port, n730_port, n731_port, n732_port, n733_port, n734_port, 
      n735_port, n736_port, n737_port, n738_port, n739_port, n740_port, 
      n741_port, n742_port, n743_port, n744_port, n745_port, n746_port, 
      n747_port, n748_port, n749_port, n750_port, n751_port, n752_port, 
      n753_port, n754_port, n755_port, n756_port, n757_port, n758_port, 
      n759_port, n760_port, n761_port, n762_port, n763_port, n764_port, 
      n765_port, n766_port, n767_port, n768_port, n769_port, n770_port, 
      n771_port, n772_port, n773_port, n774_port, n775_port, n776_port, 
      n777_port, n778_port, n779_port, n780_port, n781_port, n782_port, 
      n783_port, n784_port, n785_port, n786_port, n787_port, n788_port, 
      n789_port, n790_port, n791_port, n792_port, n793_port, n794_port, 
      n795_port, n796_port, n797_port, n798_port, n799_port, n800_port, 
      n801_port, n802_port, n803_port, n804_port, n805_port, n806_port, 
      n807_port, n808_port, n809_port, n810_port, n811_port, n812_port, 
      n813_port, n814_port, n815_port, n816_port, n817_port, n818_port, 
      n819_port, n820_port, n821_port, n822_port, n823_port, n824_port, 
      n825_port, n826_port, n827_port, n828_port, n829_port, n830_port, 
      n831_port, n832_port, n833_port, n834_port, n835_port, n836_port, 
      n837_port, n838_port, n839_port, n840_port, n841_port, n842_port, 
      n843_port, n844_port, n845_port, n846_port, n847_port, n848_port, 
      n849_port, n850_port, n851_port, n852_port, n853_port, n854_port, 
      n855_port, n856_port, n857_port, n858_port, n859_port, n860_port, 
      n861_port, n862_port, n863_port, n864_port, n865_port, n866_port, 
      n867_port, n868_port, n869_port, n870_port, n871_port, n872_port, 
      n873_port, n874_port, n875_port, n876_port, n877_port, n878_port, 
      n879_port, n880_port, n881_port, n882_port, n883_port, n884_port, 
      n885_port, n886_port, n887_port, n888_port, n889_port, n890_port, 
      n891_port, n892_port, n893_port, n894_port, n895_port, n896_port, 
      n897_port, n898_port, n899_port, n900_port, n901_port, n902_port, 
      n903_port, n904_port, n905_port, n906_port, n907_port, n908_port, 
      n909_port, n910_port, n911_port, n912_port, n913_port, n914_port, 
      n915_port, n916_port, n917_port, n918_port, n919_port, n920_port, 
      n921_port, n922_port, n923_port, n924_port, n925_port, n926_port, 
      n927_port, n928_port, n929_port, n930_port, n931_port, n932_port, 
      n933_port, n934_port, n935_port, n936_port, n937_port, n938_port, 
      n939_port, n940_port, n941_port, n942_port, n943_port, n944_port, 
      n945_port, n946_port, n947_port, n948_port, n949_port, n950_port, 
      n951_port, n952_port, n953_port, n954_port, n955_port, n956_port, 
      n957_port, n958_port, n959_port, n960_port, n961_port, n962_port, 
      n963_port, n964_port, n965_port, n966_port, n967_port, n968_port, 
      n969_port, n970_port, n971_port, n972_port, n973_port, n974_port, 
      n975_port, n976_port, n977_port, n978_port, n979_port, n980_port, 
      n981_port, n982_port, n983_port, n984_port, n985_port, n986_port, 
      n987_port, n988_port, n989_port, n990_port, n991_port, n992_port, 
      n993_port, n994_port, n995_port, n996_port, n997_port, n998_port, 
      n999_port, n1000_port, n1001_port, n1002_port, n1003_port, n1004_port, 
      n1005_port, n1006_port, n1007_port, n1008_port, n1009_port, n1010_port, 
      n1011_port, n1012_port, n1013_port, n1014_port, n1015_port, n1016_port, 
      n1017_port, n1018_port, n1019_port, n1020_port, n1021_port, n1022_port, 
      n1023_port, n1024_port, n1025_port, n1026_port, n1027_port, n1028_port, 
      n1029_port, n1030_port, n1031_port, n1032_port, n1033_port, n1034_port, 
      n1035_port, n1036_port, n1037_port, n1038_port, n1039_port, n1040_port, 
      n1041_port, n1042_port, n1043_port, n1044_port, n1045_port, n1046_port, 
      n1047_port, n1048_port, n1049_port, n1050_port, n1051_port, n1052_port, 
      n1053_port, n1054_port, n1055_port, n1056_port, n1057_port, n1058_port, 
      n1059_port, n1060_port, n1061_port, n1062_port, n1063_port, n1064_port, 
      n1065_port, n1066_port, n1067_port, n1068_port, n1069_port, n1070_port, 
      n1071_port, n1072_port, n1073_port, n1074_port, n1075_port, n1076_port, 
      n1077_port, n1078_port, n1079_port, n1080_port, n1081_port, n1082_port, 
      n1083_port, n1084_port, n1085_port, n1086_port, n1087_port, n1088_port, 
      n1089_port, n1090_port, n1091_port, n1092_port, n1093_port, n1094_port, 
      n1095_port, n1096_port, n1097_port, n1098_port, n1099_port, n1100_port, 
      n1101_port, n1102_port, n1103_port, n1104_port, n1105_port, n1106_port, 
      n1107_port, n1108_port, n1109_port, n1110_port, n1111_port, n1112_port, 
      n1113_port, n1114_port, n1115_port, n1116_port, n1117_port, n1118_port, 
      n1119_port, n1120_port, n1121_port, n1122_port, n1123_port, n1124_port, 
      n1125_port, n1126_port, n1127_port, n1128_port, n1129_port, n1130_port, 
      n1131_port, n1132_port, n1133_port, n1134_port, n1135_port, n1136_port, 
      n1137_port, n1138_port, n1139_port, n1140_port, n1141_port, n1142_port, 
      n1143_port, n1144_port, n1145_port, n1146_port, n1147_port, n1148_port, 
      n1149_port, n1150_port, n1151_port, n1152_port, n1153_port, n1154_port, 
      n1155_port, n1156_port, n1157_port, n1158_port, n1159_port, n1160_port, 
      n1161_port, n1162_port, n1163_port, n1164_port, n1165_port, n1166_port, 
      n1167_port, n1168_port, n1169_port, n1170_port, n1171_port, n1172_port, 
      n1173_port, n1174_port, n1175_port, n1176_port, n1177_port, n1178_port, 
      n1179_port, n1180_port, n1181_port, n1182_port, n1183_port, n1184_port, 
      n1185_port, n1186_port, n1187_port, n1188_port, n1189_port, n1190_port, 
      n1191_port, n1192_port, n1193_port, n1194_port, n1195_port, n1196_port, 
      n1197_port, n1198_port, n1199_port, n1200_port, n1201_port, n1202_port, 
      n1203_port, n1204_port, n1205_port, n1206_port, n1207_port, n1208_port, 
      n1209_port, n1210_port, n1211_port, n1212_port, n1213_port, n1214_port, 
      n1215_port, n1216_port, n1217_port, n1218_port, n1219_port, n1220_port, 
      n1221_port, n1222_port, n1223_port, n1224_port, n1225_port, n1226_port, 
      n1227_port, n1228_port, n1229_port, n1230_port, n1231_port, n1232_port, 
      n1233_port, n1234_port, n1235_port, n1236_port, n1237_port, n1238_port, 
      n1239_port, n1240_port, n1241_port, n1242_port, n1243_port, n1244_port, 
      n1245_port, n1246_port, n1247_port, n1248_port, n1249_port, n1250_port, 
      n1251_port, n1252_port, n1253_port, n1254_port, n1255_port, n1256_port, 
      n1257_port, n1258_port, n1259_port, n1260_port, n1261_port, n1262_port, 
      n1263_port, n1264_port, n1265_port, n1266_port, n1267_port, n1268_port, 
      n1269_port, n1270_port, n1271_port, n1272_port, n1273_port, n1274_port, 
      n1275_port, n1276_port, n1277_port, n1278_port, n1279_port, n1280_port, 
      n1281_port, n1282_port, n1283_port, n1284_port, n1285_port, n1286_port, 
      n1287_port, n1288_port, n1289_port, n1290_port, n1291_port, n1292_port, 
      n1293_port, n1294_port, n1295_port, n1296_port, n1297_port, n1298_port, 
      n1299_port, n1300_port, n1301_port, n1302_port, n1303_port, n1304_port, 
      n1305_port, n1306_port, n1307_port, n1308_port, n1309_port, n1310_port, 
      n1311_port, n1312_port, n1313_port, n1314_port, n1315_port, n1316_port, 
      n1317_port, n1318_port, n1319_port, n1320_port, n1321_port, n1322_port, 
      n1323_port, n1324_port, n1325_port, n1326_port, n1327_port, n1328_port, 
      n1329_port, n1330_port, n1331_port, n1332_port, n1333_port, n1334_port, 
      n1335_port, n1336_port, n1337_port, n1338_port, n1339_port, n1340_port, 
      n1341_port, n1342_port, n1343_port, n1344_port, n1345_port, n1346_port, 
      n1347_port, n1348_port, n1349_port, n1350_port, n1351_port, n1352_port, 
      n1353_port, n1354_port, n1355_port, n1356_port, n1357_port, n1358_port, 
      n1359_port, n1360_port, n1361_port, n1362_port, n1363_port, n1364_port, 
      n1365_port, n1366_port, n1367_port, n1368_port, n1369_port, n1370_port, 
      n1371_port, n1372_port, n1373_port, n1374_port, n1375_port, n1376_port, 
      n1377_port, n1378_port, n1379_port, n1380_port, n1381_port, n1382_port, 
      n1383_port, n1384_port, n1385_port, n1386_port, n1387_port, n1388_port, 
      n1389_port, n1390_port, n1391_port, n1392_port, n1393_port, n1394_port, 
      n1395_port, n1396_port, n1397_port, n1398_port, n1399_port, n1400_port, 
      n1401_port, n1402_port, n1403_port, n1404_port, n1405_port, n1406_port, 
      n1407_port, n1408_port, n1409_port, n1410_port, n1411_port, n1412_port, 
      n1413_port, n1414_port, n1415_port, n1416_port, n1417_port, n1418_port, 
      n1419_port, n1420_port, n1421_port, n1422_port, n1423_port, n1424_port, 
      n1425_port, n1426_port, n1427_port, n1428_port, n1429_port, n1430_port, 
      n1431_port, n1432_port, n1433_port, n1434_port, n1435_port, n1436_port, 
      n1437_port, n1438_port, n1439_port, n1440_port, n1441_port, n1442_port, 
      n1443_port, n1444_port, n1445_port, n1446_port, n1447_port, n1448_port, 
      n1449_port, n1450_port, n1451_port, n1452_port, n1453_port, n1454_port, 
      n1455_port, n1456_port, n1457_port, n1458_port, n1459_port, n1460_port, 
      n1461_port, n1462_port, n1463_port, n1464_port, n1465_port, n1466_port, 
      n1467_port, n1468_port, n1469_port, n1470_port, n1471_port, n1472_port, 
      n1473_port, n1474_port, n1475_port, n1476_port, n1477_port, n1478_port, 
      n1479_port, n1480_port, n1481_port, n1482_port, n1483_port, n1484_port, 
      n1485_port, n1486_port, n1487_port, n1488_port, n1489_port, n1490_port, 
      n1491_port, n1492_port, n1493_port, n1494_port, n1495_port, n1496_port, 
      n1497_port, n1498_port, n1499_port, n1500_port, n1501_port, n1502_port, 
      n1503_port, n1504_port, n1505_port, n1506_port, n1507_port, n1508_port, 
      n1509_port, n1510_port, n1511_port, n1512_port, n1513_port, n1514_port, 
      n1515_port, n1516_port, n1517_port, n1518_port, n1519_port, n1520_port, 
      n1521_port, n1522_port, n1523_port, n1524_port, n1525_port, n1526_port, 
      n1527_port, n1528_port, n1529_port, n1530_port, n1531_port, n1532_port, 
      n1533_port, n1534_port, n1535_port, n1536_port, n1537_port, n1538_port, 
      n1539_port, n1540_port, n1541_port, n1542_port, n1543_port, n1544_port, 
      n1545_port, n1546_port, n1547_port, n1548_port, n1549_port, n1550_port, 
      n1551_port, n1552_port, n1553_port, n1554_port, n1555_port, n1556_port, 
      n1557_port, n1558_port, n1559_port, n1560_port, n1561_port, n1562_port, 
      n1563_port, n1564_port, n1565_port, n1566_port, n1567_port, n1568_port, 
      n1569_port, n1570_port, n1571_port, n1572_port, n1573_port, n1574_port, 
      n1575_port, n1576_port, n1577_port, n1578_port, n1579_port, n1580_port, 
      n1581_port, n1582_port, n1583_port, n1584_port, n1585_port, n1586_port, 
      n1587_port, n1588_port, n1589_port, n1590_port, n1591_port, n1592_port, 
      n1593_port, n1594_port, n1595_port, n1596_port, n1597_port, n1598_port, 
      n1599_port, n1600_port, n1601_port, n1602_port, n1603_port, n1604_port, 
      n1605_port, n1606_port, n1607_port, n1608_port, n1609_port, n1610_port, 
      n1611_port, n1612_port, n1613_port, n1614_port, n1615_port, n1616_port, 
      n1617_port, n1618_port, n1619_port, n1620_port, n1621_port, n1622_port, 
      n1623_port, n1624_port, n1625_port, n1626_port, n1627_port, n1628_port, 
      n1629_port, n1630_port, n1631_port, n1632_port, n1633_port, n1634_port, 
      n1635_port, n1636_port, n1637_port, n1638_port, n1639_port, n1640_port, 
      n1641_port, n1642_port, n1643_port, n1644_port, n1645_port, n1646_port, 
      n1647_port, n1648_port, n1649_port, n1650_port, n1651_port, n1652_port, 
      n1653_port, n1654_port, n1655_port, n1656_port, n1657_port, n1658_port, 
      n1659_port, n1660_port, n1661_port, n1662_port, n1663_port, n1664_port, 
      n1665_port, n1666_port, n1667_port, n1668_port, n1669_port, n1670_port, 
      n1671_port, n1672_port, n1673_port, n1674_port, n1675_port, n1676_port, 
      n1677_port, n1678_port, n1679_port, n1680_port, n1681_port, n1682_port, 
      n1683_port, n1684_port, n1685_port, n1686_port, n1687_port, n1688_port, 
      n1689_port, n1690_port, n1691_port, n1692_port, n1693_port, n1694_port, 
      n1695_port, n1696_port, n1697_port, n1698_port, n1699_port, n1700_port, 
      n1701_port, n1702_port, n1703_port, n1704_port, n1705_port, n1706_port, 
      n1707_port, n1708_port, n1709_port, n1710_port, n1711_port, n1712_port, 
      n1713_port, n1714_port, n1715_port, n1716_port, n1717_port, n1718_port, 
      n1719_port, n1720_port, n1721_port, n1722_port, n1723_port, n1724_port, 
      n1725_port, n1726_port, n1727_port, n1728_port, n1729_port, n1730_port, 
      n1731_port, n1732_port, n1733_port, n1734_port, n1735_port, n1736_port, 
      n1737_port, n1738_port, n1739_port, n1740_port, n1741_port, n1742_port, 
      n1743_port, n1744_port, n1745_port, n1746_port, n1747_port, n1748_port, 
      n1749_port, n1750_port, n1751_port, n1752_port, n1753_port, n1754_port, 
      n1755_port, n1756_port, n1757_port, n1758_port, n1759_port, n1760_port, 
      n1761_port, n1762_port, n1763_port, n1764_port, n1765_port, n1766_port, 
      n1767_port, n1768_port, n1769_port, n1770_port, n1771_port, n1772_port, 
      n1773_port, n1774_port, n1775_port, n1776_port, n1777_port, n1778_port, 
      n1779_port, n1780_port, n1781_port, n1782_port, n1783_port, n1784_port, 
      n1785_port, n1786_port, n1787_port, n1788_port, n1789_port, n1790_port, 
      n1791_port, n1792_port, n1793_port, n1794_port, n1795_port, n1796_port, 
      n1797_port, n1798_port, n1799_port, n1800_port, n1801_port, n1802_port, 
      n1803_port, n1804_port, n1805_port, n1806_port, n1807_port, n1808_port, 
      n1809_port, n1810_port, n1811_port, n1812_port, n1813_port, n1814_port, 
      n1815_port, n1816_port, n1817_port, n1818_port, n1819_port, n1820_port, 
      n1821_port, n1822_port, n1823_port, n1824_port, n1825_port, n1826_port, 
      n1827_port, n1828_port, n1829_port, n1830_port, n1831_port, n1832_port, 
      n1833_port, n1834_port, n1835_port, n1836_port, n1837_port, n1838_port, 
      n1839_port, n1840_port, n1841_port, n1842_port, n1843_port, n1844_port, 
      n1845_port, n1846_port, n1847_port, n1848_port, n1849_port, n1850_port, 
      n1851_port, n1852_port, n1853_port, n1854_port, n1855_port, n1856_port, 
      n1857_port, n1858_port, n1859_port, n1860_port, n1861_port, n1862_port, 
      n1863_port, n1864_port, n1865_port, n1866_port, n1867_port, n1868_port, 
      n1869_port, n1870_port, n1871_port, n1872_port, n1873_port, n1874_port, 
      n1875_port, n1876_port, n1877_port, n1878_port, n1879_port, n1880_port, 
      n1881_port, n1882_port, n1883_port, n1884_port, n1885_port, n1886_port, 
      n1887_port, n1888_port, n1889_port, n1890_port, n1891_port, n1892_port, 
      n1893_port, n1894_port, n1895_port, n1896_port, n1897_port, n1898_port, 
      n1899_port, n1900_port, n1901_port, n1902_port, n1903_port, n1904_port, 
      n1905_port, n1906_port, n1907_port, n1908_port, n1909_port, n1910_port, 
      n1911_port, n1912_port, n1913_port, n1914_port, n1915_port, n1916_port, 
      n1917_port, n1918_port, n1919_port, n1920_port, n1921_port, n1922_port, 
      n1923_port, n1924_port, n1925_port, n1926_port, n1927_port, n1928_port, 
      n1929_port, n1930_port, n1931_port, n1932_port, n1933_port, n1934_port, 
      n1935_port, n1936_port, n1937_port, n1938_port, n1939_port, n1940_port, 
      n1941_port, n1942_port, n1943_port, n1944_port, n1945_port, n1946_port, 
      n1947_port, n1948_port, n1949_port, n1950_port, n1951_port, n1952_port, 
      n1953_port, n1954_port, n1955_port, n1956_port, n1957_port, n1958_port, 
      n1959_port, n1960_port, n1961_port, n1962_port, n1963_port, n1964_port, 
      n1965_port, n1966_port, n1967_port, n1968_port, n1969_port, n1970_port, 
      n1971_port, n1972_port, n1973_port, n1974_port, n1975_port, n1976_port, 
      n1977_port, n1978_port, n1979_port, n1980_port, n1981_port, n1982_port, 
      n1983_port, n1984_port, n1985_port, n1986_port, n1987_port, n1988_port, 
      n1989_port, n1990_port, n1991_port, n1992_port, n1993_port, n1994_port, 
      n1995_port, n1996_port, n1997_port, n1998_port, n1999_port, n2000_port, 
      n2001_port, n2002_port, n2003_port, n2004_port, n2005_port, n2006_port, 
      n2007_port, n2008_port, n2009_port, n2010_port, n2011_port, n2012_port, 
      n2013_port, n2014_port, n2015_port, n2016_port, n2017_port, n2018_port, 
      n2019_port, n2020_port, n2021_port, n2022_port, n2023_port, n2024_port, 
      n2025_port, n2026_port, n2027_port, n2028_port, n2029_port, n2030_port, 
      n2031_port, n2032_port, n2033_port, n2034_port, n2035_port, n2036_port, 
      n2037_port, n2038_port, n2039_port, n2040_port, n2041_port, n2042_port, 
      n2043_port, n2044_port, n2045_port, n2046_port, n2047_port, n2048_port, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
      n6246, n6247, n6248, n6249, n7211, n7212, n7213, n7214, n7215, n7216, 
      n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, 
      n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, 
      n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, 
      n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, 
      n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, 
      n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, 
      n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, 
      n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, 
      n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, 
      n7307, n7308, n7309, n7310, n7311, n7312, n7318, n7319, n7320, n7321, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8498, 
      n8499, n8500, n8501, n8504, n8505, n8506, n8507, n8508, n8509, n8510, 
      n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, 
      n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, 
      n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, 
      n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, 
      n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, 
      n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, 
      n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, 
      n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, 
      n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, 
      n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, 
      n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, 
      n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, 
      n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, 
      n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, 
      n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, 
      n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, 
      n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, 
      n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, 
      n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, 
      n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, 
      n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, 
      n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, 
      n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, 
      n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, 
      n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, 
      n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, 
      n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, 
      n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, 
      n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, 
      n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, 
      n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, 
      n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, 
      n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, 
      n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, 
      n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, 
      n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, 
      n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, 
      n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, 
      n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, 
      n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, 
      n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, 
      n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, 
      n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, 
      n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, 
      n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, 
      n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, 
      n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, 
      n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, 
      n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, 
      n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, 
      n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, 
      n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, 
      n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, 
      n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, 
      n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, 
      n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, 
      n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, 
      n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, 
      n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, 
      n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, 
      n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, 
      n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, 
      n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, 
      n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, 
      n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, 
      n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, 
      n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, 
      n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, 
      n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, 
      n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, 
      n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, 
      n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, 
      n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
      n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, 
      n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, 
      n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, 
      n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, 
      n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, 
      n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, 
      n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, 
      n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, 
      n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, 
      n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, 
      n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, 
      n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, 
      n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, 
      n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, 
      n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, 
      n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, 
      n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, 
      n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, 
      n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, 
      n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, 
      n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, 
      n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, 
      n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, 
      n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, 
      n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, 
      n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, 
      n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, 
      n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, 
      n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, 
      n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, 
      n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, 
      n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, 
      n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, 
      n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, 
      n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, 
      n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, 
      n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, 
      n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, 
      n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, 
      n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, 
      n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, 
      n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
      n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, 
      n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, 
      n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, 
      n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, 
      n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, 
      n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, 
      n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, 
      n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, 
      n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, 
      n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, 
      n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, 
      n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, 
      n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, 
      n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, 
      n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, 
      n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, 
      n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, 
      n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, 
      n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, 
      n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, 
      n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, 
      n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, 
      n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, 
      n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, 
      n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, 
      n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, 
      n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, 
      n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, 
      n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, 
      n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
      n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, 
      n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, 
      n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, 
      n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, 
      n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, 
      n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, 
      n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
      n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, 
      n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, 
      n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, 
      n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, 
      n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, 
      n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, 
      n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, 
      n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, 
      n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, 
      n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, 
      n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, 
      n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, 
      n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, 
      n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, 
      n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, 
      n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, 
      n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, 
      n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, 
      n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, 
      n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, 
      n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
      n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, 
      n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, 
      n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, 
      n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, 
      n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, 
      n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, 
      n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, 
      n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, 
      n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, 
      n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, 
      n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, 
      n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, 
      n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, 
      n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, 
      n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, 
      n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, 
      n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, 
      n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, 
      n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, 
      n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, 
      n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, 
      n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, 
      n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, 
      n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, 
      n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, 
      n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, 
      n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, 
      n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, 
      n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, 
      n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, 
      n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, 
      n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, 
      n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, 
      n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, 
      n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, 
      n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, 
      n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, 
      n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, 
      n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, 
      n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
      n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, 
      n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, 
      n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, 
      n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, 
      n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, 
      n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, 
      n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, 
      n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, 
      n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, 
      n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, 
      n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, 
      n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, 
      n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, 
      n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, 
      n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, 
      n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, 
      n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, 
      n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, 
      n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, 
      n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, 
      n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, 
      n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, 
      n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, 
      n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, 
      n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, 
      n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, 
      n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, 
      n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, 
      n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, 
      n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, 
      n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, 
      n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, 
      n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, 
      n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, 
      n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, 
      n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, 
      n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, 
      n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, 
      n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, 
      n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, 
      n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, 
      n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, 
      n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, 
      n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, 
      n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, 
      n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, 
      n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, 
      n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, 
      n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, 
      n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, 
      n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, 
      n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, 
      n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, 
      n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, 
      n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, 
      n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, 
      n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, 
      n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, 
      n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, 
      n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, 
      n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, 
      n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, 
      n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, 
      n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, 
      n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, 
      n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, 
      n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, 
      n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, 
      n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, 
      n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, 
      n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, 
      n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, 
      n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, 
      n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
      n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, 
      n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, 
      n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, 
      n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, 
      n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, 
      n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, 
      n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, 
      n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, 
      n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, 
      n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, 
      n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, 
      n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, 
      n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, 
      n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, 
      n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, 
      n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, 
      n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, 
      n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, 
      n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, 
      n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, 
      n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, 
      n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, 
      n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, 
      n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, 
      n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, 
      n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, 
      n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, 
      n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
      n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, 
      n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, 
      n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, 
      n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, 
      n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, 
      n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, 
      n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, 
      n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, 
      n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, 
      n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, 
      n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, 
      n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, 
      n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, 
      n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, 
      n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, 
      n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, 
      n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, 
      n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, 
      n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, 
      n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, 
      n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, 
      n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, 
      n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, 
      n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, 
      n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, 
      n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, 
      n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, 
      n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, 
      n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, 
      n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, 
      n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, 
      n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, 
      n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, 
      n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, 
      n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, 
      n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, 
      n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, 
      n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, 
      n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, 
      n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, 
      n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, 
      n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, 
      n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, 
      n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, 
      n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, 
      n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, 
      n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, 
      n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, 
      n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, 
      n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, 
      n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, 
      n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, 
      n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, 
      n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, 
      n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, 
      n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, 
      n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, 
      n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, 
      n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, 
      n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, 
      n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, 
      n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, 
      n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, 
      n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, 
      n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, 
      n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, 
      n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, 
      n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, 
      n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, 
      n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, 
      n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, 
      n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, 
      n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, 
      n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, 
      n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, 
      n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, 
      n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, 
      n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, 
      n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, 
      n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, 
      n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, 
      n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, 
      n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, 
      n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, 
      n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, 
      n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, 
      n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, 
      n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, 
      n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, 
      n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, 
      n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, 
      n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, 
      n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, 
      n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, 
      n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, 
      n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, 
      n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, 
      n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, 
      n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, 
      n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, 
      n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, 
      n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, 
      n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, 
      n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, 
      n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, 
      n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, 
      n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, 
      n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, 
      n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, 
      n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, 
      n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, 
      n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, 
      n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, 
      n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, 
      n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, 
      n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, 
      n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, 
      n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, 
      n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, 
      n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, 
      n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, 
      n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, 
      n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, 
      n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, 
      n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, 
      n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, 
      n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, 
      n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, 
      n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, 
      n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, 
      n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, 
      n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087 : std_logic;

begin
   
   OUT1_reg_63_inst : DLH_X1 port map( G => n12184, D => N2071, Q => OUT1(63));
   OUT1_reg_62_inst : DLH_X1 port map( G => n12184, D => N2072, Q => OUT1(62));
   OUT1_reg_61_inst : DLH_X1 port map( G => n12184, D => N2073, Q => OUT1(61));
   OUT1_reg_60_inst : DLH_X1 port map( G => n12184, D => N2074, Q => OUT1(60));
   OUT1_reg_59_inst : DLH_X1 port map( G => n12184, D => N2075, Q => OUT1(59));
   OUT1_reg_58_inst : DLH_X1 port map( G => n12184, D => N2076, Q => OUT1(58));
   OUT1_reg_57_inst : DLH_X1 port map( G => n12184, D => N2077, Q => OUT1(57));
   OUT1_reg_56_inst : DLH_X1 port map( G => n12184, D => N2078, Q => OUT1(56));
   OUT1_reg_55_inst : DLH_X1 port map( G => n12184, D => N2079, Q => OUT1(55));
   OUT1_reg_54_inst : DLH_X1 port map( G => n12183, D => N2080, Q => OUT1(54));
   OUT1_reg_53_inst : DLH_X1 port map( G => n12183, D => N2081, Q => OUT1(53));
   OUT1_reg_52_inst : DLH_X1 port map( G => n12183, D => N2082, Q => OUT1(52));
   OUT1_reg_51_inst : DLH_X1 port map( G => n12183, D => N2083, Q => OUT1(51));
   OUT1_reg_50_inst : DLH_X1 port map( G => n12183, D => N2084, Q => OUT1(50));
   OUT1_reg_49_inst : DLH_X1 port map( G => n12183, D => N2085, Q => OUT1(49));
   OUT1_reg_48_inst : DLH_X1 port map( G => n12183, D => N2086, Q => OUT1(48));
   OUT1_reg_47_inst : DLH_X1 port map( G => n12183, D => N2087, Q => OUT1(47));
   OUT1_reg_46_inst : DLH_X1 port map( G => n12183, D => N2088, Q => OUT1(46));
   OUT1_reg_45_inst : DLH_X1 port map( G => n12183, D => N2089, Q => OUT1(45));
   OUT1_reg_44_inst : DLH_X1 port map( G => n12183, D => N2090, Q => OUT1(44));
   OUT1_reg_43_inst : DLH_X1 port map( G => n12182, D => N2091, Q => OUT1(43));
   OUT1_reg_42_inst : DLH_X1 port map( G => n12182, D => N2092, Q => OUT1(42));
   OUT1_reg_41_inst : DLH_X1 port map( G => n12182, D => N2093, Q => OUT1(41));
   OUT1_reg_40_inst : DLH_X1 port map( G => n12182, D => N2094, Q => OUT1(40));
   OUT1_reg_39_inst : DLH_X1 port map( G => n12182, D => N2095, Q => OUT1(39));
   OUT1_reg_38_inst : DLH_X1 port map( G => n12182, D => N2096, Q => OUT1(38));
   OUT1_reg_37_inst : DLH_X1 port map( G => n12182, D => N2097, Q => OUT1(37));
   OUT1_reg_36_inst : DLH_X1 port map( G => n12182, D => N2098, Q => OUT1(36));
   OUT1_reg_35_inst : DLH_X1 port map( G => n12182, D => N2099, Q => OUT1(35));
   OUT1_reg_34_inst : DLH_X1 port map( G => n12182, D => N2100, Q => OUT1(34));
   OUT1_reg_33_inst : DLH_X1 port map( G => n12182, D => N2101, Q => OUT1(33));
   OUT1_reg_32_inst : DLH_X1 port map( G => n12181, D => N2102, Q => OUT1(32));
   OUT1_reg_31_inst : DLH_X1 port map( G => n12181, D => N2103, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => n12181, D => N2104, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => n12181, D => N2105, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => n12181, D => N2106, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => n12181, D => N2107, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => n12181, D => N2108, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => n12181, D => N2109, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => n12181, D => N2110, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => n12181, D => N2111, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => n12181, D => N2112, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => n12180, D => N2113, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => n12180, D => N2114, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => n12180, D => N2115, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => n12180, D => N2116, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => n12180, D => N2117, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => n12180, D => N2118, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => n12180, D => N2119, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => n12180, D => N2120, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => n12180, D => N2121, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => n12180, D => N2122, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => n12180, D => N2123, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => n12179, D => N2124, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => n12179, D => N2125, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => n12179, D => N2126, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => n12179, D => N2127, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => n12179, D => N2128, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => n12179, D => N2129, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => n12179, D => N2130, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => n12179, D => N2131, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => n12179, D => N2132, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => n12179, D => N2133, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => n12179, D => N2134, Q => OUT1(0));
   OUT2_reg_63_inst : DLH_X1 port map( G => n12176, D => N2136, Q => OUT2(63));
   OUT2_reg_62_inst : DLH_X1 port map( G => n12176, D => N2137, Q => OUT2(62));
   OUT2_reg_61_inst : DLH_X1 port map( G => n12176, D => N2138, Q => OUT2(61));
   OUT2_reg_60_inst : DLH_X1 port map( G => n12176, D => N2139, Q => OUT2(60));
   OUT2_reg_59_inst : DLH_X1 port map( G => n12176, D => N2140, Q => OUT2(59));
   OUT2_reg_58_inst : DLH_X1 port map( G => n12176, D => N2141, Q => OUT2(58));
   OUT2_reg_57_inst : DLH_X1 port map( G => n12176, D => N2142, Q => OUT2(57));
   OUT2_reg_56_inst : DLH_X1 port map( G => n12176, D => N2143, Q => OUT2(56));
   OUT2_reg_55_inst : DLH_X1 port map( G => n12176, D => N2144, Q => OUT2(55));
   OUT2_reg_54_inst : DLH_X1 port map( G => n12175, D => N2145, Q => OUT2(54));
   OUT2_reg_53_inst : DLH_X1 port map( G => n12175, D => N2146, Q => OUT2(53));
   OUT2_reg_52_inst : DLH_X1 port map( G => n12175, D => N2147, Q => OUT2(52));
   OUT2_reg_51_inst : DLH_X1 port map( G => n12175, D => N2148, Q => OUT2(51));
   OUT2_reg_50_inst : DLH_X1 port map( G => n12175, D => N2149, Q => OUT2(50));
   OUT2_reg_49_inst : DLH_X1 port map( G => n12175, D => N2150, Q => OUT2(49));
   OUT2_reg_48_inst : DLH_X1 port map( G => n12175, D => N2151, Q => OUT2(48));
   OUT2_reg_47_inst : DLH_X1 port map( G => n12175, D => N2152, Q => OUT2(47));
   OUT2_reg_46_inst : DLH_X1 port map( G => n12175, D => N2153, Q => OUT2(46));
   OUT2_reg_45_inst : DLH_X1 port map( G => n12175, D => N2154, Q => OUT2(45));
   OUT2_reg_44_inst : DLH_X1 port map( G => n12175, D => N2155, Q => OUT2(44));
   OUT2_reg_43_inst : DLH_X1 port map( G => n12174, D => N2156, Q => OUT2(43));
   OUT2_reg_42_inst : DLH_X1 port map( G => n12174, D => N2157, Q => OUT2(42));
   OUT2_reg_41_inst : DLH_X1 port map( G => n12174, D => N2158, Q => OUT2(41));
   OUT2_reg_40_inst : DLH_X1 port map( G => n12174, D => N2159, Q => OUT2(40));
   OUT2_reg_39_inst : DLH_X1 port map( G => n12174, D => N2160, Q => OUT2(39));
   OUT2_reg_38_inst : DLH_X1 port map( G => n12174, D => N2161, Q => OUT2(38));
   OUT2_reg_37_inst : DLH_X1 port map( G => n12174, D => N2162, Q => OUT2(37));
   OUT2_reg_36_inst : DLH_X1 port map( G => n12174, D => N2163, Q => OUT2(36));
   OUT2_reg_35_inst : DLH_X1 port map( G => n12174, D => N2164, Q => OUT2(35));
   OUT2_reg_34_inst : DLH_X1 port map( G => n12174, D => N2165, Q => OUT2(34));
   OUT2_reg_33_inst : DLH_X1 port map( G => n12174, D => N2166, Q => OUT2(33));
   OUT2_reg_32_inst : DLH_X1 port map( G => n12173, D => N2167, Q => OUT2(32));
   OUT2_reg_31_inst : DLH_X1 port map( G => n12173, D => N2168, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n12173, D => N2169, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n12173, D => N2170, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n12173, D => N2171, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n12173, D => N2172, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n12173, D => N2173, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n12173, D => N2174, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n12173, D => N2175, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n12173, D => N2176, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n12173, D => N2177, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n12172, D => N2178, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n12172, D => N2179, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n12172, D => N2180, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n12172, D => N2181, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n12172, D => N2182, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n12172, D => N2183, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n12172, D => N2184, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n12172, D => N2185, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n12172, D => N2186, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n12172, D => N2187, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n12172, D => N2188, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n12171, D => N2189, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n12171, D => N2190, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n12171, D => N2191, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n12171, D => N2192, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n12171, D => N2193, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n12171, D => N2194, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n12171, D => N2195, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n12171, D => N2196, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n12171, D => N2197, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n12171, D => N2198, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n12171, D => N2199, Q => OUT2(0));
   NEXT_REGISTERS_reg_0_63_inst : DLH_X1 port map( G => n11883, D => N4313, Q 
                           => NEXT_REGISTERS_0_63_port);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => N2069, CK => CLK, Q => n9966
                           , QN => n1);
   NEXT_REGISTERS_reg_0_62_inst : DLH_X1 port map( G => n11883, D => N4312, Q 
                           => NEXT_REGISTERS_0_62_port);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => N2068, CK => CLK, Q => n9964
                           , QN => n2);
   NEXT_REGISTERS_reg_0_61_inst : DLH_X1 port map( G => n11883, D => N4311, Q 
                           => NEXT_REGISTERS_0_61_port);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => N2067, CK => CLK, Q => n9962
                           , QN => n3);
   NEXT_REGISTERS_reg_0_60_inst : DLH_X1 port map( G => n11883, D => N4310, Q 
                           => NEXT_REGISTERS_0_60_port);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => N2066, CK => CLK, Q => n9960
                           , QN => n4);
   NEXT_REGISTERS_reg_0_59_inst : DLH_X1 port map( G => n11883, D => N4309, Q 
                           => NEXT_REGISTERS_0_59_port);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => N2065, CK => CLK, Q => n9958
                           , QN => n5);
   NEXT_REGISTERS_reg_0_58_inst : DLH_X1 port map( G => n11883, D => N4308, Q 
                           => NEXT_REGISTERS_0_58_port);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => N2064, CK => CLK, Q => n9956
                           , QN => n6);
   NEXT_REGISTERS_reg_0_57_inst : DLH_X1 port map( G => n11883, D => N4307, Q 
                           => NEXT_REGISTERS_0_57_port);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => N2063, CK => CLK, Q => n9954
                           , QN => n7);
   NEXT_REGISTERS_reg_0_56_inst : DLH_X1 port map( G => n11883, D => N4306, Q 
                           => NEXT_REGISTERS_0_56_port);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => N2062, CK => CLK, Q => n9952
                           , QN => n8);
   NEXT_REGISTERS_reg_0_55_inst : DLH_X1 port map( G => n11883, D => N4305, Q 
                           => NEXT_REGISTERS_0_55_port);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => N2061, CK => CLK, Q => n9950
                           , QN => n9);
   NEXT_REGISTERS_reg_0_54_inst : DLH_X1 port map( G => n11883, D => N4304, Q 
                           => NEXT_REGISTERS_0_54_port);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => N2060, CK => CLK, Q => n9948
                           , QN => n10);
   NEXT_REGISTERS_reg_0_53_inst : DLH_X1 port map( G => n11883, D => N4303, Q 
                           => NEXT_REGISTERS_0_53_port);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => N2059, CK => CLK, Q => n9946
                           , QN => n11);
   NEXT_REGISTERS_reg_0_52_inst : DLH_X1 port map( G => n11884, D => N4302, Q 
                           => NEXT_REGISTERS_0_52_port);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => N2058, CK => CLK, Q => n9944
                           , QN => n12);
   NEXT_REGISTERS_reg_0_51_inst : DLH_X1 port map( G => n11884, D => N4301, Q 
                           => NEXT_REGISTERS_0_51_port);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => N2057, CK => CLK, Q => n9942
                           , QN => n13);
   NEXT_REGISTERS_reg_0_50_inst : DLH_X1 port map( G => n11884, D => N4300, Q 
                           => NEXT_REGISTERS_0_50_port);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => N2056, CK => CLK, Q => n9940
                           , QN => n14);
   NEXT_REGISTERS_reg_0_49_inst : DLH_X1 port map( G => n11884, D => N4299, Q 
                           => NEXT_REGISTERS_0_49_port);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => N2055, CK => CLK, Q => n9938
                           , QN => n15);
   NEXT_REGISTERS_reg_0_48_inst : DLH_X1 port map( G => n11884, D => N4298, Q 
                           => NEXT_REGISTERS_0_48_port);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => N2054, CK => CLK, Q => n9936
                           , QN => n16);
   NEXT_REGISTERS_reg_0_47_inst : DLH_X1 port map( G => n11884, D => N4297, Q 
                           => NEXT_REGISTERS_0_47_port);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => N2053, CK => CLK, Q => n9934
                           , QN => n17);
   NEXT_REGISTERS_reg_0_46_inst : DLH_X1 port map( G => n11884, D => N4296, Q 
                           => NEXT_REGISTERS_0_46_port);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => N2052, CK => CLK, Q => n9932
                           , QN => n18);
   NEXT_REGISTERS_reg_0_45_inst : DLH_X1 port map( G => n11884, D => N4295, Q 
                           => NEXT_REGISTERS_0_45_port);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => N2051, CK => CLK, Q => n9930
                           , QN => n19);
   NEXT_REGISTERS_reg_0_44_inst : DLH_X1 port map( G => n11884, D => N4294, Q 
                           => NEXT_REGISTERS_0_44_port);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => N2050, CK => CLK, Q => n9928
                           , QN => n20);
   NEXT_REGISTERS_reg_0_43_inst : DLH_X1 port map( G => n11884, D => N4293, Q 
                           => NEXT_REGISTERS_0_43_port);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => N2049, CK => CLK, Q => n9926
                           , QN => n21);
   NEXT_REGISTERS_reg_0_42_inst : DLH_X1 port map( G => n11884, D => N4292, Q 
                           => NEXT_REGISTERS_0_42_port);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => N2048, CK => CLK, Q => n9924
                           , QN => n22_port);
   NEXT_REGISTERS_reg_0_41_inst : DLH_X1 port map( G => n11885, D => N4291, Q 
                           => NEXT_REGISTERS_0_41_port);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => N2047, CK => CLK, Q => n9922
                           , QN => n23_port);
   NEXT_REGISTERS_reg_0_40_inst : DLH_X1 port map( G => n11885, D => N4290, Q 
                           => NEXT_REGISTERS_0_40_port);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => N2046, CK => CLK, Q => n9920
                           , QN => n24_port);
   NEXT_REGISTERS_reg_0_39_inst : DLH_X1 port map( G => n11885, D => N4289, Q 
                           => NEXT_REGISTERS_0_39_port);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => N2045, CK => CLK, Q => n9918
                           , QN => n25_port);
   NEXT_REGISTERS_reg_0_38_inst : DLH_X1 port map( G => n11885, D => N4288, Q 
                           => NEXT_REGISTERS_0_38_port);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => N2044, CK => CLK, Q => n9916
                           , QN => n26_port);
   NEXT_REGISTERS_reg_0_37_inst : DLH_X1 port map( G => n11885, D => N4287, Q 
                           => NEXT_REGISTERS_0_37_port);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => N2043, CK => CLK, Q => n9914
                           , QN => n27_port);
   NEXT_REGISTERS_reg_0_36_inst : DLH_X1 port map( G => n11885, D => N4286, Q 
                           => NEXT_REGISTERS_0_36_port);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => N2042, CK => CLK, Q => n9912
                           , QN => n28_port);
   NEXT_REGISTERS_reg_0_35_inst : DLH_X1 port map( G => n11885, D => N4285, Q 
                           => NEXT_REGISTERS_0_35_port);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => N2041, CK => CLK, Q => n9910
                           , QN => n29_port);
   NEXT_REGISTERS_reg_0_34_inst : DLH_X1 port map( G => n11885, D => N4284, Q 
                           => NEXT_REGISTERS_0_34_port);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => N2040, CK => CLK, Q => n9908
                           , QN => n30_port);
   NEXT_REGISTERS_reg_0_33_inst : DLH_X1 port map( G => n11885, D => N4283, Q 
                           => NEXT_REGISTERS_0_33_port);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => N2039, CK => CLK, Q => n9906
                           , QN => n31_port);
   NEXT_REGISTERS_reg_0_32_inst : DLH_X1 port map( G => n11885, D => N4282, Q 
                           => NEXT_REGISTERS_0_32_port);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => N2038, CK => CLK, Q => n9904
                           , QN => n32_port);
   NEXT_REGISTERS_reg_0_31_inst : DLH_X1 port map( G => n11885, D => N4281, Q 
                           => NEXT_REGISTERS_0_31_port);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => N2037, CK => CLK, Q => n9902
                           , QN => n33_port);
   NEXT_REGISTERS_reg_0_30_inst : DLH_X1 port map( G => n11886, D => N4280, Q 
                           => NEXT_REGISTERS_0_30_port);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => N2036, CK => CLK, Q => n9900
                           , QN => n34_port);
   NEXT_REGISTERS_reg_0_29_inst : DLH_X1 port map( G => n11886, D => N4279, Q 
                           => NEXT_REGISTERS_0_29_port);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => N2035, CK => CLK, Q => n9898
                           , QN => n35_port);
   NEXT_REGISTERS_reg_0_28_inst : DLH_X1 port map( G => n11886, D => N4278, Q 
                           => NEXT_REGISTERS_0_28_port);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => N2034, CK => CLK, Q => n9896
                           , QN => n36_port);
   NEXT_REGISTERS_reg_0_27_inst : DLH_X1 port map( G => n11886, D => N4277, Q 
                           => NEXT_REGISTERS_0_27_port);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => N2033, CK => CLK, Q => n9894
                           , QN => n37_port);
   NEXT_REGISTERS_reg_0_26_inst : DLH_X1 port map( G => n11886, D => N4276, Q 
                           => NEXT_REGISTERS_0_26_port);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => N2032, CK => CLK, Q => n9892
                           , QN => n38_port);
   NEXT_REGISTERS_reg_0_25_inst : DLH_X1 port map( G => n11886, D => N4275, Q 
                           => NEXT_REGISTERS_0_25_port);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => N2031, CK => CLK, Q => n9890
                           , QN => n39_port);
   NEXT_REGISTERS_reg_0_24_inst : DLH_X1 port map( G => n11886, D => N4274, Q 
                           => NEXT_REGISTERS_0_24_port);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => N2030, CK => CLK, Q => n9888
                           , QN => n40_port);
   NEXT_REGISTERS_reg_0_23_inst : DLH_X1 port map( G => n11886, D => N4273, Q 
                           => NEXT_REGISTERS_0_23_port);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => N2029, CK => CLK, Q => n9886
                           , QN => n41_port);
   NEXT_REGISTERS_reg_0_22_inst : DLH_X1 port map( G => n11886, D => N4272, Q 
                           => NEXT_REGISTERS_0_22_port);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => N2028, CK => CLK, Q => n9884
                           , QN => n42_port);
   NEXT_REGISTERS_reg_0_21_inst : DLH_X1 port map( G => n11886, D => N4271, Q 
                           => NEXT_REGISTERS_0_21_port);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => N2027, CK => CLK, Q => n9882
                           , QN => n43_port);
   NEXT_REGISTERS_reg_0_20_inst : DLH_X1 port map( G => n11886, D => N4270, Q 
                           => NEXT_REGISTERS_0_20_port);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => N2026, CK => CLK, Q => n9880
                           , QN => n44_port);
   NEXT_REGISTERS_reg_0_19_inst : DLH_X1 port map( G => n11887, D => N4269, Q 
                           => NEXT_REGISTERS_0_19_port);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => N2025, CK => CLK, Q => n9878
                           , QN => n45_port);
   NEXT_REGISTERS_reg_0_18_inst : DLH_X1 port map( G => n11887, D => N4268, Q 
                           => NEXT_REGISTERS_0_18_port);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => N2024, CK => CLK, Q => n9876
                           , QN => n46_port);
   NEXT_REGISTERS_reg_0_17_inst : DLH_X1 port map( G => n11887, D => N4267, Q 
                           => NEXT_REGISTERS_0_17_port);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => N2023, CK => CLK, Q => n9874
                           , QN => n47_port);
   NEXT_REGISTERS_reg_0_16_inst : DLH_X1 port map( G => n11887, D => N4266, Q 
                           => NEXT_REGISTERS_0_16_port);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => N2022, CK => CLK, Q => n9872
                           , QN => n48_port);
   NEXT_REGISTERS_reg_0_15_inst : DLH_X1 port map( G => n11887, D => N4265, Q 
                           => NEXT_REGISTERS_0_15_port);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => N2021, CK => CLK, Q => n9870
                           , QN => n49_port);
   NEXT_REGISTERS_reg_0_14_inst : DLH_X1 port map( G => n11887, D => N4264, Q 
                           => NEXT_REGISTERS_0_14_port);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => N2020, CK => CLK, Q => n9868
                           , QN => n50_port);
   NEXT_REGISTERS_reg_0_13_inst : DLH_X1 port map( G => n11887, D => N4263, Q 
                           => NEXT_REGISTERS_0_13_port);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => N2019, CK => CLK, Q => n9866
                           , QN => n51_port);
   NEXT_REGISTERS_reg_0_12_inst : DLH_X1 port map( G => n11887, D => N4262, Q 
                           => NEXT_REGISTERS_0_12_port);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => N2018, CK => CLK, Q => n9864
                           , QN => n52_port);
   NEXT_REGISTERS_reg_0_11_inst : DLH_X1 port map( G => n11887, D => N4261, Q 
                           => NEXT_REGISTERS_0_11_port);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => N2017, CK => CLK, Q => n9862
                           , QN => n53_port);
   NEXT_REGISTERS_reg_0_10_inst : DLH_X1 port map( G => n11887, D => N4260, Q 
                           => NEXT_REGISTERS_0_10_port);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => N2016, CK => CLK, Q => n9860
                           , QN => n54_port);
   NEXT_REGISTERS_reg_0_9_inst : DLH_X1 port map( G => n11887, D => N4259, Q =>
                           NEXT_REGISTERS_0_9_port);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => N2015, CK => CLK, Q => n9858,
                           QN => n55_port);
   NEXT_REGISTERS_reg_0_8_inst : DLH_X1 port map( G => n11888, D => N4258, Q =>
                           NEXT_REGISTERS_0_8_port);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => N2014, CK => CLK, Q => n9856,
                           QN => n56_port);
   NEXT_REGISTERS_reg_0_7_inst : DLH_X1 port map( G => n11888, D => N4257, Q =>
                           NEXT_REGISTERS_0_7_port);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => N2013, CK => CLK, Q => n9854,
                           QN => n57_port);
   NEXT_REGISTERS_reg_0_6_inst : DLH_X1 port map( G => n11888, D => N4256, Q =>
                           NEXT_REGISTERS_0_6_port);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => N2012, CK => CLK, Q => n9852,
                           QN => n58_port);
   NEXT_REGISTERS_reg_0_5_inst : DLH_X1 port map( G => n11888, D => N4255, Q =>
                           NEXT_REGISTERS_0_5_port);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => N2011, CK => CLK, Q => n9850,
                           QN => n59_port);
   NEXT_REGISTERS_reg_0_4_inst : DLH_X1 port map( G => n11888, D => N4254, Q =>
                           NEXT_REGISTERS_0_4_port);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => N2010, CK => CLK, Q => n9848,
                           QN => n60_port);
   NEXT_REGISTERS_reg_0_3_inst : DLH_X1 port map( G => n11888, D => N4253, Q =>
                           NEXT_REGISTERS_0_3_port);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => N2009, CK => CLK, Q => n9846,
                           QN => n61_port);
   NEXT_REGISTERS_reg_0_2_inst : DLH_X1 port map( G => n11888, D => N4252, Q =>
                           NEXT_REGISTERS_0_2_port);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => N2008, CK => CLK, Q => n9844,
                           QN => n62_port);
   NEXT_REGISTERS_reg_0_1_inst : DLH_X1 port map( G => n11888, D => N4251, Q =>
                           NEXT_REGISTERS_0_1_port);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => N2007, CK => CLK, Q => n9842,
                           QN => n63_port);
   NEXT_REGISTERS_reg_0_0_inst : DLH_X1 port map( G => n11888, D => N4250, Q =>
                           NEXT_REGISTERS_0_0_port);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => N2006, CK => CLK, Q => n9840,
                           QN => n64_port);
   NEXT_REGISTERS_reg_1_63_inst : DLH_X1 port map( G => n11892, D => N4248, Q 
                           => NEXT_REGISTERS_1_63_port);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => N2005, CK => CLK, Q => 
                           n_1000, QN => n65_port);
   NEXT_REGISTERS_reg_1_62_inst : DLH_X1 port map( G => n11892, D => N4247, Q 
                           => NEXT_REGISTERS_1_62_port);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => N2004, CK => CLK, Q => 
                           n_1001, QN => n66_port);
   NEXT_REGISTERS_reg_1_61_inst : DLH_X1 port map( G => n11892, D => N4246, Q 
                           => NEXT_REGISTERS_1_61_port);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => N2003, CK => CLK, Q => 
                           n_1002, QN => n67_port);
   NEXT_REGISTERS_reg_1_60_inst : DLH_X1 port map( G => n11892, D => N4245, Q 
                           => NEXT_REGISTERS_1_60_port);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => N2002, CK => CLK, Q => 
                           n_1003, QN => n68_port);
   NEXT_REGISTERS_reg_1_59_inst : DLH_X1 port map( G => n11892, D => N4244, Q 
                           => NEXT_REGISTERS_1_59_port);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => N2001, CK => CLK, Q => 
                           n_1004, QN => n69_port);
   NEXT_REGISTERS_reg_1_58_inst : DLH_X1 port map( G => n11892, D => N4243, Q 
                           => NEXT_REGISTERS_1_58_port);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => N2000, CK => CLK, Q => 
                           n_1005, QN => n70_port);
   NEXT_REGISTERS_reg_1_57_inst : DLH_X1 port map( G => n11892, D => N4242, Q 
                           => NEXT_REGISTERS_1_57_port);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => N1999, CK => CLK, Q => 
                           n_1006, QN => n71_port);
   NEXT_REGISTERS_reg_1_56_inst : DLH_X1 port map( G => n11892, D => N4241, Q 
                           => NEXT_REGISTERS_1_56_port);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => N1998, CK => CLK, Q => 
                           n_1007, QN => n72_port);
   NEXT_REGISTERS_reg_1_55_inst : DLH_X1 port map( G => n11892, D => N4240, Q 
                           => NEXT_REGISTERS_1_55_port);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => N1997, CK => CLK, Q => 
                           n_1008, QN => n73_port);
   NEXT_REGISTERS_reg_1_54_inst : DLH_X1 port map( G => n11892, D => N4239, Q 
                           => NEXT_REGISTERS_1_54_port);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => N1996, CK => CLK, Q => 
                           n_1009, QN => n74_port);
   NEXT_REGISTERS_reg_1_53_inst : DLH_X1 port map( G => n11892, D => N4238, Q 
                           => NEXT_REGISTERS_1_53_port);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => N1995, CK => CLK, Q => 
                           n_1010, QN => n75_port);
   NEXT_REGISTERS_reg_1_52_inst : DLH_X1 port map( G => n11893, D => N4237, Q 
                           => NEXT_REGISTERS_1_52_port);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => N1994, CK => CLK, Q => 
                           n_1011, QN => n76_port);
   NEXT_REGISTERS_reg_1_51_inst : DLH_X1 port map( G => n11893, D => N4236, Q 
                           => NEXT_REGISTERS_1_51_port);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => N1993, CK => CLK, Q => 
                           n_1012, QN => n77_port);
   NEXT_REGISTERS_reg_1_50_inst : DLH_X1 port map( G => n11893, D => N4235, Q 
                           => NEXT_REGISTERS_1_50_port);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => N1992, CK => CLK, Q => 
                           n_1013, QN => n78_port);
   NEXT_REGISTERS_reg_1_49_inst : DLH_X1 port map( G => n11893, D => N4234, Q 
                           => NEXT_REGISTERS_1_49_port);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => N1991, CK => CLK, Q => 
                           n_1014, QN => n79_port);
   NEXT_REGISTERS_reg_1_48_inst : DLH_X1 port map( G => n11893, D => N4233, Q 
                           => NEXT_REGISTERS_1_48_port);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => N1990, CK => CLK, Q => 
                           n_1015, QN => n80_port);
   NEXT_REGISTERS_reg_1_47_inst : DLH_X1 port map( G => n11893, D => N4232, Q 
                           => NEXT_REGISTERS_1_47_port);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => N1989, CK => CLK, Q => 
                           n_1016, QN => n81_port);
   NEXT_REGISTERS_reg_1_46_inst : DLH_X1 port map( G => n11893, D => N4231, Q 
                           => NEXT_REGISTERS_1_46_port);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => N1988, CK => CLK, Q => 
                           n_1017, QN => n82_port);
   NEXT_REGISTERS_reg_1_45_inst : DLH_X1 port map( G => n11893, D => N4230, Q 
                           => NEXT_REGISTERS_1_45_port);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => N1987, CK => CLK, Q => 
                           n_1018, QN => n83_port);
   NEXT_REGISTERS_reg_1_44_inst : DLH_X1 port map( G => n11893, D => N4229, Q 
                           => NEXT_REGISTERS_1_44_port);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => N1986, CK => CLK, Q => 
                           n_1019, QN => n84_port);
   NEXT_REGISTERS_reg_1_43_inst : DLH_X1 port map( G => n11893, D => N4228, Q 
                           => NEXT_REGISTERS_1_43_port);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => N1985, CK => CLK, Q => 
                           n_1020, QN => n85_port);
   NEXT_REGISTERS_reg_1_42_inst : DLH_X1 port map( G => n11893, D => N4227, Q 
                           => NEXT_REGISTERS_1_42_port);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => N1984, CK => CLK, Q => 
                           n_1021, QN => n86_port);
   NEXT_REGISTERS_reg_1_41_inst : DLH_X1 port map( G => n11894, D => N4226, Q 
                           => NEXT_REGISTERS_1_41_port);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => N1983, CK => CLK, Q => 
                           n_1022, QN => n87_port);
   NEXT_REGISTERS_reg_1_40_inst : DLH_X1 port map( G => n11894, D => N4225, Q 
                           => NEXT_REGISTERS_1_40_port);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => N1982, CK => CLK, Q => 
                           n_1023, QN => n88_port);
   NEXT_REGISTERS_reg_1_39_inst : DLH_X1 port map( G => n11894, D => N4224, Q 
                           => NEXT_REGISTERS_1_39_port);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => N1981, CK => CLK, Q => 
                           n_1024, QN => n89_port);
   NEXT_REGISTERS_reg_1_38_inst : DLH_X1 port map( G => n11894, D => N4223, Q 
                           => NEXT_REGISTERS_1_38_port);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => N1980, CK => CLK, Q => 
                           n_1025, QN => n90_port);
   NEXT_REGISTERS_reg_1_37_inst : DLH_X1 port map( G => n11894, D => N4222, Q 
                           => NEXT_REGISTERS_1_37_port);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => N1979, CK => CLK, Q => 
                           n_1026, QN => n91_port);
   NEXT_REGISTERS_reg_1_36_inst : DLH_X1 port map( G => n11894, D => N4221, Q 
                           => NEXT_REGISTERS_1_36_port);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => N1978, CK => CLK, Q => 
                           n_1027, QN => n92_port);
   NEXT_REGISTERS_reg_1_35_inst : DLH_X1 port map( G => n11894, D => N4220, Q 
                           => NEXT_REGISTERS_1_35_port);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => N1977, CK => CLK, Q => 
                           n_1028, QN => n93_port);
   NEXT_REGISTERS_reg_1_34_inst : DLH_X1 port map( G => n11894, D => N4219, Q 
                           => NEXT_REGISTERS_1_34_port);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => N1976, CK => CLK, Q => 
                           n_1029, QN => n94_port);
   NEXT_REGISTERS_reg_1_33_inst : DLH_X1 port map( G => n11894, D => N4218, Q 
                           => NEXT_REGISTERS_1_33_port);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => N1975, CK => CLK, Q => 
                           n_1030, QN => n95_port);
   NEXT_REGISTERS_reg_1_32_inst : DLH_X1 port map( G => n11894, D => N4217, Q 
                           => NEXT_REGISTERS_1_32_port);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => N1974, CK => CLK, Q => 
                           n_1031, QN => n96_port);
   NEXT_REGISTERS_reg_1_31_inst : DLH_X1 port map( G => n11894, D => N4216, Q 
                           => NEXT_REGISTERS_1_31_port);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => N1973, CK => CLK, Q => 
                           n_1032, QN => n97_port);
   NEXT_REGISTERS_reg_1_30_inst : DLH_X1 port map( G => n11895, D => N4215, Q 
                           => NEXT_REGISTERS_1_30_port);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => N1972, CK => CLK, Q => 
                           n_1033, QN => n98_port);
   NEXT_REGISTERS_reg_1_29_inst : DLH_X1 port map( G => n11895, D => N4214, Q 
                           => NEXT_REGISTERS_1_29_port);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => N1971, CK => CLK, Q => 
                           n_1034, QN => n99_port);
   NEXT_REGISTERS_reg_1_28_inst : DLH_X1 port map( G => n11895, D => N4213, Q 
                           => NEXT_REGISTERS_1_28_port);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => N1970, CK => CLK, Q => 
                           n_1035, QN => n100_port);
   NEXT_REGISTERS_reg_1_27_inst : DLH_X1 port map( G => n11895, D => N4212, Q 
                           => NEXT_REGISTERS_1_27_port);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => N1969, CK => CLK, Q => 
                           n_1036, QN => n101_port);
   NEXT_REGISTERS_reg_1_26_inst : DLH_X1 port map( G => n11895, D => N4211, Q 
                           => NEXT_REGISTERS_1_26_port);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => N1968, CK => CLK, Q => 
                           n_1037, QN => n102_port);
   NEXT_REGISTERS_reg_1_25_inst : DLH_X1 port map( G => n11895, D => N4210, Q 
                           => NEXT_REGISTERS_1_25_port);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => N1967, CK => CLK, Q => 
                           n_1038, QN => n103_port);
   NEXT_REGISTERS_reg_1_24_inst : DLH_X1 port map( G => n11895, D => N4209, Q 
                           => NEXT_REGISTERS_1_24_port);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => N1966, CK => CLK, Q => 
                           n_1039, QN => n104_port);
   NEXT_REGISTERS_reg_1_23_inst : DLH_X1 port map( G => n11895, D => N4208, Q 
                           => NEXT_REGISTERS_1_23_port);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => N1965, CK => CLK, Q => 
                           n_1040, QN => n105_port);
   NEXT_REGISTERS_reg_1_22_inst : DLH_X1 port map( G => n11895, D => N4207, Q 
                           => NEXT_REGISTERS_1_22_port);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => N1964, CK => CLK, Q => 
                           n_1041, QN => n106_port);
   NEXT_REGISTERS_reg_1_21_inst : DLH_X1 port map( G => n11895, D => N4206, Q 
                           => NEXT_REGISTERS_1_21_port);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => N1963, CK => CLK, Q => 
                           n_1042, QN => n107_port);
   NEXT_REGISTERS_reg_1_20_inst : DLH_X1 port map( G => n11895, D => N4205, Q 
                           => NEXT_REGISTERS_1_20_port);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => N1962, CK => CLK, Q => 
                           n_1043, QN => n108_port);
   NEXT_REGISTERS_reg_1_19_inst : DLH_X1 port map( G => n11896, D => N4204, Q 
                           => NEXT_REGISTERS_1_19_port);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => N1961, CK => CLK, Q => 
                           n_1044, QN => n109_port);
   NEXT_REGISTERS_reg_1_18_inst : DLH_X1 port map( G => n11896, D => N4203, Q 
                           => NEXT_REGISTERS_1_18_port);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => N1960, CK => CLK, Q => 
                           n_1045, QN => n110_port);
   NEXT_REGISTERS_reg_1_17_inst : DLH_X1 port map( G => n11896, D => N4202, Q 
                           => NEXT_REGISTERS_1_17_port);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => N1959, CK => CLK, Q => 
                           n_1046, QN => n111_port);
   NEXT_REGISTERS_reg_1_16_inst : DLH_X1 port map( G => n11896, D => N4201, Q 
                           => NEXT_REGISTERS_1_16_port);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => N1958, CK => CLK, Q => 
                           n_1047, QN => n112_port);
   NEXT_REGISTERS_reg_1_15_inst : DLH_X1 port map( G => n11896, D => N4200, Q 
                           => NEXT_REGISTERS_1_15_port);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => N1957, CK => CLK, Q => 
                           n_1048, QN => n113_port);
   NEXT_REGISTERS_reg_1_14_inst : DLH_X1 port map( G => n11896, D => N4199, Q 
                           => NEXT_REGISTERS_1_14_port);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => N1956, CK => CLK, Q => 
                           n_1049, QN => n114_port);
   NEXT_REGISTERS_reg_1_13_inst : DLH_X1 port map( G => n11896, D => N4198, Q 
                           => NEXT_REGISTERS_1_13_port);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => N1955, CK => CLK, Q => 
                           n_1050, QN => n115_port);
   NEXT_REGISTERS_reg_1_12_inst : DLH_X1 port map( G => n11896, D => N4197, Q 
                           => NEXT_REGISTERS_1_12_port);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => N1954, CK => CLK, Q => 
                           n_1051, QN => n116_port);
   NEXT_REGISTERS_reg_1_11_inst : DLH_X1 port map( G => n11896, D => N4196, Q 
                           => NEXT_REGISTERS_1_11_port);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => N1953, CK => CLK, Q => 
                           n_1052, QN => n117_port);
   NEXT_REGISTERS_reg_1_10_inst : DLH_X1 port map( G => n11896, D => N4195, Q 
                           => NEXT_REGISTERS_1_10_port);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => N1952, CK => CLK, Q => 
                           n_1053, QN => n118_port);
   NEXT_REGISTERS_reg_1_9_inst : DLH_X1 port map( G => n11896, D => N4194, Q =>
                           NEXT_REGISTERS_1_9_port);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => N1951, CK => CLK, Q => n_1054
                           , QN => n119_port);
   NEXT_REGISTERS_reg_1_8_inst : DLH_X1 port map( G => n11897, D => N4193, Q =>
                           NEXT_REGISTERS_1_8_port);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => N1950, CK => CLK, Q => n_1055
                           , QN => n120_port);
   NEXT_REGISTERS_reg_1_7_inst : DLH_X1 port map( G => n11897, D => N4192, Q =>
                           NEXT_REGISTERS_1_7_port);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => N1949, CK => CLK, Q => n_1056
                           , QN => n121_port);
   NEXT_REGISTERS_reg_1_6_inst : DLH_X1 port map( G => n11897, D => N4191, Q =>
                           NEXT_REGISTERS_1_6_port);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => N1948, CK => CLK, Q => n_1057
                           , QN => n122_port);
   NEXT_REGISTERS_reg_1_5_inst : DLH_X1 port map( G => n11897, D => N4190, Q =>
                           NEXT_REGISTERS_1_5_port);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => N1947, CK => CLK, Q => n_1058
                           , QN => n123_port);
   NEXT_REGISTERS_reg_1_4_inst : DLH_X1 port map( G => n11897, D => N4189, Q =>
                           NEXT_REGISTERS_1_4_port);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => N1946, CK => CLK, Q => n_1059
                           , QN => n124_port);
   NEXT_REGISTERS_reg_1_3_inst : DLH_X1 port map( G => n11897, D => N4188, Q =>
                           NEXT_REGISTERS_1_3_port);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => N1945, CK => CLK, Q => n_1060
                           , QN => n125_port);
   NEXT_REGISTERS_reg_1_2_inst : DLH_X1 port map( G => n11897, D => N4187, Q =>
                           NEXT_REGISTERS_1_2_port);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => N1944, CK => CLK, Q => n_1061
                           , QN => n126_port);
   NEXT_REGISTERS_reg_1_1_inst : DLH_X1 port map( G => n11897, D => N4186, Q =>
                           NEXT_REGISTERS_1_1_port);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => N1943, CK => CLK, Q => n_1062
                           , QN => n127_port);
   NEXT_REGISTERS_reg_1_0_inst : DLH_X1 port map( G => n11897, D => N4185, Q =>
                           NEXT_REGISTERS_1_0_port);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => N1942, CK => CLK, Q => n_1063
                           , QN => n128_port);
   NEXT_REGISTERS_reg_2_63_inst : DLH_X1 port map( G => n11901, D => N4183, Q 
                           => NEXT_REGISTERS_2_63_port);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => N1941, CK => CLK, Q => 
                           n10414, QN => n129_port);
   NEXT_REGISTERS_reg_2_62_inst : DLH_X1 port map( G => n11901, D => N4182, Q 
                           => NEXT_REGISTERS_2_62_port);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => N1940, CK => CLK, Q => 
                           n10412, QN => n130_port);
   NEXT_REGISTERS_reg_2_61_inst : DLH_X1 port map( G => n11901, D => N4181, Q 
                           => NEXT_REGISTERS_2_61_port);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => N1939, CK => CLK, Q => 
                           n10410, QN => n131_port);
   NEXT_REGISTERS_reg_2_60_inst : DLH_X1 port map( G => n11901, D => N4180, Q 
                           => NEXT_REGISTERS_2_60_port);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => N1938, CK => CLK, Q => 
                           n10408, QN => n132_port);
   NEXT_REGISTERS_reg_2_59_inst : DLH_X1 port map( G => n11901, D => N4179, Q 
                           => NEXT_REGISTERS_2_59_port);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => N1937, CK => CLK, Q => 
                           n10406, QN => n133_port);
   NEXT_REGISTERS_reg_2_58_inst : DLH_X1 port map( G => n11901, D => N4178, Q 
                           => NEXT_REGISTERS_2_58_port);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => N1936, CK => CLK, Q => 
                           n10404, QN => n134_port);
   NEXT_REGISTERS_reg_2_57_inst : DLH_X1 port map( G => n11901, D => N4177, Q 
                           => NEXT_REGISTERS_2_57_port);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => N1935, CK => CLK, Q => 
                           n10402, QN => n135_port);
   NEXT_REGISTERS_reg_2_56_inst : DLH_X1 port map( G => n11901, D => N4176, Q 
                           => NEXT_REGISTERS_2_56_port);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => N1934, CK => CLK, Q => 
                           n10400, QN => n136_port);
   NEXT_REGISTERS_reg_2_55_inst : DLH_X1 port map( G => n11901, D => N4175, Q 
                           => NEXT_REGISTERS_2_55_port);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => N1933, CK => CLK, Q => 
                           n10398, QN => n137_port);
   NEXT_REGISTERS_reg_2_54_inst : DLH_X1 port map( G => n11901, D => N4174, Q 
                           => NEXT_REGISTERS_2_54_port);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => N1932, CK => CLK, Q => 
                           n10396, QN => n138_port);
   NEXT_REGISTERS_reg_2_53_inst : DLH_X1 port map( G => n11901, D => N4173, Q 
                           => NEXT_REGISTERS_2_53_port);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => N1931, CK => CLK, Q => 
                           n10394, QN => n139_port);
   NEXT_REGISTERS_reg_2_52_inst : DLH_X1 port map( G => n11902, D => N4172, Q 
                           => NEXT_REGISTERS_2_52_port);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => N1930, CK => CLK, Q => 
                           n10392, QN => n140_port);
   NEXT_REGISTERS_reg_2_51_inst : DLH_X1 port map( G => n11902, D => N4171, Q 
                           => NEXT_REGISTERS_2_51_port);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => N1929, CK => CLK, Q => 
                           n10390, QN => n141_port);
   NEXT_REGISTERS_reg_2_50_inst : DLH_X1 port map( G => n11902, D => N4170, Q 
                           => NEXT_REGISTERS_2_50_port);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => N1928, CK => CLK, Q => 
                           n10388, QN => n142_port);
   NEXT_REGISTERS_reg_2_49_inst : DLH_X1 port map( G => n11902, D => N4169, Q 
                           => NEXT_REGISTERS_2_49_port);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => N1927, CK => CLK, Q => 
                           n10386, QN => n143_port);
   NEXT_REGISTERS_reg_2_48_inst : DLH_X1 port map( G => n11902, D => N4168, Q 
                           => NEXT_REGISTERS_2_48_port);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => N1926, CK => CLK, Q => 
                           n10384, QN => n144_port);
   NEXT_REGISTERS_reg_2_47_inst : DLH_X1 port map( G => n11902, D => N4167, Q 
                           => NEXT_REGISTERS_2_47_port);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => N1925, CK => CLK, Q => 
                           n10382, QN => n145_port);
   NEXT_REGISTERS_reg_2_46_inst : DLH_X1 port map( G => n11902, D => N4166, Q 
                           => NEXT_REGISTERS_2_46_port);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => N1924, CK => CLK, Q => 
                           n10380, QN => n146_port);
   NEXT_REGISTERS_reg_2_45_inst : DLH_X1 port map( G => n11902, D => N4165, Q 
                           => NEXT_REGISTERS_2_45_port);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => N1923, CK => CLK, Q => 
                           n10378, QN => n147_port);
   NEXT_REGISTERS_reg_2_44_inst : DLH_X1 port map( G => n11902, D => N4164, Q 
                           => NEXT_REGISTERS_2_44_port);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => N1922, CK => CLK, Q => 
                           n10376, QN => n148_port);
   NEXT_REGISTERS_reg_2_43_inst : DLH_X1 port map( G => n11902, D => N4163, Q 
                           => NEXT_REGISTERS_2_43_port);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => N1921, CK => CLK, Q => 
                           n10374, QN => n149_port);
   NEXT_REGISTERS_reg_2_42_inst : DLH_X1 port map( G => n11902, D => N4162, Q 
                           => NEXT_REGISTERS_2_42_port);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => N1920, CK => CLK, Q => 
                           n10372, QN => n150_port);
   NEXT_REGISTERS_reg_2_41_inst : DLH_X1 port map( G => n11903, D => N4161, Q 
                           => NEXT_REGISTERS_2_41_port);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => N1919, CK => CLK, Q => 
                           n10370, QN => n151_port);
   NEXT_REGISTERS_reg_2_40_inst : DLH_X1 port map( G => n11903, D => N4160, Q 
                           => NEXT_REGISTERS_2_40_port);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => N1918, CK => CLK, Q => 
                           n10368, QN => n152_port);
   NEXT_REGISTERS_reg_2_39_inst : DLH_X1 port map( G => n11903, D => N4159, Q 
                           => NEXT_REGISTERS_2_39_port);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => N1917, CK => CLK, Q => 
                           n10366, QN => n153_port);
   NEXT_REGISTERS_reg_2_38_inst : DLH_X1 port map( G => n11903, D => N4158, Q 
                           => NEXT_REGISTERS_2_38_port);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => N1916, CK => CLK, Q => 
                           n10364, QN => n154_port);
   NEXT_REGISTERS_reg_2_37_inst : DLH_X1 port map( G => n11903, D => N4157, Q 
                           => NEXT_REGISTERS_2_37_port);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => N1915, CK => CLK, Q => 
                           n10362, QN => n155_port);
   NEXT_REGISTERS_reg_2_36_inst : DLH_X1 port map( G => n11903, D => N4156, Q 
                           => NEXT_REGISTERS_2_36_port);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => N1914, CK => CLK, Q => 
                           n10360, QN => n156_port);
   NEXT_REGISTERS_reg_2_35_inst : DLH_X1 port map( G => n11903, D => N4155, Q 
                           => NEXT_REGISTERS_2_35_port);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => N1913, CK => CLK, Q => 
                           n10358, QN => n157_port);
   NEXT_REGISTERS_reg_2_34_inst : DLH_X1 port map( G => n11903, D => N4154, Q 
                           => NEXT_REGISTERS_2_34_port);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => N1912, CK => CLK, Q => 
                           n10356, QN => n158_port);
   NEXT_REGISTERS_reg_2_33_inst : DLH_X1 port map( G => n11903, D => N4153, Q 
                           => NEXT_REGISTERS_2_33_port);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => N1911, CK => CLK, Q => 
                           n10354, QN => n159_port);
   NEXT_REGISTERS_reg_2_32_inst : DLH_X1 port map( G => n11903, D => N4152, Q 
                           => NEXT_REGISTERS_2_32_port);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => N1910, CK => CLK, Q => 
                           n10352, QN => n160_port);
   NEXT_REGISTERS_reg_2_31_inst : DLH_X1 port map( G => n11903, D => N4151, Q 
                           => NEXT_REGISTERS_2_31_port);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => N1909, CK => CLK, Q => 
                           n10350, QN => n161_port);
   NEXT_REGISTERS_reg_2_30_inst : DLH_X1 port map( G => n11904, D => N4150, Q 
                           => NEXT_REGISTERS_2_30_port);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => N1908, CK => CLK, Q => 
                           n10348, QN => n162_port);
   NEXT_REGISTERS_reg_2_29_inst : DLH_X1 port map( G => n11904, D => N4149, Q 
                           => NEXT_REGISTERS_2_29_port);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => N1907, CK => CLK, Q => 
                           n10346, QN => n163_port);
   NEXT_REGISTERS_reg_2_28_inst : DLH_X1 port map( G => n11904, D => N4148, Q 
                           => NEXT_REGISTERS_2_28_port);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => N1906, CK => CLK, Q => 
                           n10344, QN => n164_port);
   NEXT_REGISTERS_reg_2_27_inst : DLH_X1 port map( G => n11904, D => N4147, Q 
                           => NEXT_REGISTERS_2_27_port);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => N1905, CK => CLK, Q => 
                           n10342, QN => n165_port);
   NEXT_REGISTERS_reg_2_26_inst : DLH_X1 port map( G => n11904, D => N4146, Q 
                           => NEXT_REGISTERS_2_26_port);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => N1904, CK => CLK, Q => 
                           n10340, QN => n166_port);
   NEXT_REGISTERS_reg_2_25_inst : DLH_X1 port map( G => n11904, D => N4145, Q 
                           => NEXT_REGISTERS_2_25_port);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => N1903, CK => CLK, Q => 
                           n10338, QN => n167_port);
   NEXT_REGISTERS_reg_2_24_inst : DLH_X1 port map( G => n11904, D => N4144, Q 
                           => NEXT_REGISTERS_2_24_port);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => N1902, CK => CLK, Q => 
                           n10336, QN => n168_port);
   NEXT_REGISTERS_reg_2_23_inst : DLH_X1 port map( G => n11904, D => N4143, Q 
                           => NEXT_REGISTERS_2_23_port);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => N1901, CK => CLK, Q => 
                           n10334, QN => n169_port);
   NEXT_REGISTERS_reg_2_22_inst : DLH_X1 port map( G => n11904, D => N4142, Q 
                           => NEXT_REGISTERS_2_22_port);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => N1900, CK => CLK, Q => 
                           n10332, QN => n170_port);
   NEXT_REGISTERS_reg_2_21_inst : DLH_X1 port map( G => n11904, D => N4141, Q 
                           => NEXT_REGISTERS_2_21_port);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => N1899, CK => CLK, Q => 
                           n10330, QN => n171_port);
   NEXT_REGISTERS_reg_2_20_inst : DLH_X1 port map( G => n11904, D => N4140, Q 
                           => NEXT_REGISTERS_2_20_port);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => N1898, CK => CLK, Q => 
                           n10328, QN => n172_port);
   NEXT_REGISTERS_reg_2_19_inst : DLH_X1 port map( G => n11905, D => N4139, Q 
                           => NEXT_REGISTERS_2_19_port);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => N1897, CK => CLK, Q => 
                           n10326, QN => n173_port);
   NEXT_REGISTERS_reg_2_18_inst : DLH_X1 port map( G => n11905, D => N4138, Q 
                           => NEXT_REGISTERS_2_18_port);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => N1896, CK => CLK, Q => 
                           n10324, QN => n174_port);
   NEXT_REGISTERS_reg_2_17_inst : DLH_X1 port map( G => n11905, D => N4137, Q 
                           => NEXT_REGISTERS_2_17_port);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => N1895, CK => CLK, Q => 
                           n10322, QN => n175_port);
   NEXT_REGISTERS_reg_2_16_inst : DLH_X1 port map( G => n11905, D => N4136, Q 
                           => NEXT_REGISTERS_2_16_port);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => N1894, CK => CLK, Q => 
                           n10320, QN => n176_port);
   NEXT_REGISTERS_reg_2_15_inst : DLH_X1 port map( G => n11905, D => N4135, Q 
                           => NEXT_REGISTERS_2_15_port);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => N1893, CK => CLK, Q => 
                           n10318, QN => n177_port);
   NEXT_REGISTERS_reg_2_14_inst : DLH_X1 port map( G => n11905, D => N4134, Q 
                           => NEXT_REGISTERS_2_14_port);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => N1892, CK => CLK, Q => 
                           n10316, QN => n178_port);
   NEXT_REGISTERS_reg_2_13_inst : DLH_X1 port map( G => n11905, D => N4133, Q 
                           => NEXT_REGISTERS_2_13_port);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => N1891, CK => CLK, Q => 
                           n10314, QN => n179_port);
   NEXT_REGISTERS_reg_2_12_inst : DLH_X1 port map( G => n11905, D => N4132, Q 
                           => NEXT_REGISTERS_2_12_port);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => N1890, CK => CLK, Q => 
                           n10312, QN => n180_port);
   NEXT_REGISTERS_reg_2_11_inst : DLH_X1 port map( G => n11905, D => N4131, Q 
                           => NEXT_REGISTERS_2_11_port);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => N1889, CK => CLK, Q => 
                           n10310, QN => n181_port);
   NEXT_REGISTERS_reg_2_10_inst : DLH_X1 port map( G => n11905, D => N4130, Q 
                           => NEXT_REGISTERS_2_10_port);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => N1888, CK => CLK, Q => 
                           n10308, QN => n182_port);
   NEXT_REGISTERS_reg_2_9_inst : DLH_X1 port map( G => n11905, D => N4129, Q =>
                           NEXT_REGISTERS_2_9_port);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => N1887, CK => CLK, Q => n10306
                           , QN => n183_port);
   NEXT_REGISTERS_reg_2_8_inst : DLH_X1 port map( G => n11906, D => N4128, Q =>
                           NEXT_REGISTERS_2_8_port);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => N1886, CK => CLK, Q => n10304
                           , QN => n184_port);
   NEXT_REGISTERS_reg_2_7_inst : DLH_X1 port map( G => n11906, D => N4127, Q =>
                           NEXT_REGISTERS_2_7_port);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => N1885, CK => CLK, Q => n10302
                           , QN => n185_port);
   NEXT_REGISTERS_reg_2_6_inst : DLH_X1 port map( G => n11906, D => N4126, Q =>
                           NEXT_REGISTERS_2_6_port);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => N1884, CK => CLK, Q => n10300
                           , QN => n186_port);
   NEXT_REGISTERS_reg_2_5_inst : DLH_X1 port map( G => n11906, D => N4125, Q =>
                           NEXT_REGISTERS_2_5_port);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => N1883, CK => CLK, Q => n10298
                           , QN => n187_port);
   NEXT_REGISTERS_reg_2_4_inst : DLH_X1 port map( G => n11906, D => N4124, Q =>
                           NEXT_REGISTERS_2_4_port);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => N1882, CK => CLK, Q => n10296
                           , QN => n188_port);
   NEXT_REGISTERS_reg_2_3_inst : DLH_X1 port map( G => n11906, D => N4123, Q =>
                           NEXT_REGISTERS_2_3_port);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => N1881, CK => CLK, Q => n10294
                           , QN => n189_port);
   NEXT_REGISTERS_reg_2_2_inst : DLH_X1 port map( G => n11906, D => N4122, Q =>
                           NEXT_REGISTERS_2_2_port);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => N1880, CK => CLK, Q => n10292
                           , QN => n190_port);
   NEXT_REGISTERS_reg_2_1_inst : DLH_X1 port map( G => n11906, D => N4121, Q =>
                           NEXT_REGISTERS_2_1_port);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => N1879, CK => CLK, Q => n10290
                           , QN => n191_port);
   NEXT_REGISTERS_reg_2_0_inst : DLH_X1 port map( G => n11906, D => N4120, Q =>
                           NEXT_REGISTERS_2_0_port);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => N1878, CK => CLK, Q => n10288
                           , QN => n192_port);
   NEXT_REGISTERS_reg_3_63_inst : DLH_X1 port map( G => n11910, D => N4118, Q 
                           => NEXT_REGISTERS_3_63_port);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => N1877, CK => CLK, Q => 
                           n_1064, QN => n193_port);
   NEXT_REGISTERS_reg_3_62_inst : DLH_X1 port map( G => n11910, D => N4117, Q 
                           => NEXT_REGISTERS_3_62_port);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => N1876, CK => CLK, Q => 
                           n_1065, QN => n194_port);
   NEXT_REGISTERS_reg_3_61_inst : DLH_X1 port map( G => n11910, D => N4116, Q 
                           => NEXT_REGISTERS_3_61_port);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => N1875, CK => CLK, Q => 
                           n_1066, QN => n195_port);
   NEXT_REGISTERS_reg_3_60_inst : DLH_X1 port map( G => n11910, D => N4115, Q 
                           => NEXT_REGISTERS_3_60_port);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => N1874, CK => CLK, Q => 
                           n_1067, QN => n196_port);
   NEXT_REGISTERS_reg_3_59_inst : DLH_X1 port map( G => n11910, D => N4114, Q 
                           => NEXT_REGISTERS_3_59_port);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => N1873, CK => CLK, Q => 
                           n_1068, QN => n197_port);
   NEXT_REGISTERS_reg_3_58_inst : DLH_X1 port map( G => n11910, D => N4113, Q 
                           => NEXT_REGISTERS_3_58_port);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => N1872, CK => CLK, Q => 
                           n_1069, QN => n198_port);
   NEXT_REGISTERS_reg_3_57_inst : DLH_X1 port map( G => n11910, D => N4112, Q 
                           => NEXT_REGISTERS_3_57_port);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => N1871, CK => CLK, Q => 
                           n_1070, QN => n199_port);
   NEXT_REGISTERS_reg_3_56_inst : DLH_X1 port map( G => n11910, D => N4111, Q 
                           => NEXT_REGISTERS_3_56_port);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => N1870, CK => CLK, Q => 
                           n_1071, QN => n200_port);
   NEXT_REGISTERS_reg_3_55_inst : DLH_X1 port map( G => n11910, D => N4110, Q 
                           => NEXT_REGISTERS_3_55_port);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => N1869, CK => CLK, Q => 
                           n_1072, QN => n201_port);
   NEXT_REGISTERS_reg_3_54_inst : DLH_X1 port map( G => n11910, D => N4109, Q 
                           => NEXT_REGISTERS_3_54_port);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => N1868, CK => CLK, Q => 
                           n_1073, QN => n202_port);
   NEXT_REGISTERS_reg_3_53_inst : DLH_X1 port map( G => n11910, D => N4108, Q 
                           => NEXT_REGISTERS_3_53_port);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => N1867, CK => CLK, Q => 
                           n_1074, QN => n203_port);
   NEXT_REGISTERS_reg_3_52_inst : DLH_X1 port map( G => n11911, D => N4107, Q 
                           => NEXT_REGISTERS_3_52_port);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => N1866, CK => CLK, Q => 
                           n_1075, QN => n204_port);
   NEXT_REGISTERS_reg_3_51_inst : DLH_X1 port map( G => n11911, D => N4106, Q 
                           => NEXT_REGISTERS_3_51_port);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => N1865, CK => CLK, Q => 
                           n_1076, QN => n205_port);
   NEXT_REGISTERS_reg_3_50_inst : DLH_X1 port map( G => n11911, D => N4105, Q 
                           => NEXT_REGISTERS_3_50_port);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => N1864, CK => CLK, Q => 
                           n_1077, QN => n206_port);
   NEXT_REGISTERS_reg_3_49_inst : DLH_X1 port map( G => n11911, D => N4104, Q 
                           => NEXT_REGISTERS_3_49_port);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => N1863, CK => CLK, Q => 
                           n_1078, QN => n207_port);
   NEXT_REGISTERS_reg_3_48_inst : DLH_X1 port map( G => n11911, D => N4103, Q 
                           => NEXT_REGISTERS_3_48_port);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => N1862, CK => CLK, Q => 
                           n_1079, QN => n208_port);
   NEXT_REGISTERS_reg_3_47_inst : DLH_X1 port map( G => n11911, D => N4102, Q 
                           => NEXT_REGISTERS_3_47_port);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => N1861, CK => CLK, Q => 
                           n_1080, QN => n209_port);
   NEXT_REGISTERS_reg_3_46_inst : DLH_X1 port map( G => n11911, D => N4101, Q 
                           => NEXT_REGISTERS_3_46_port);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => N1860, CK => CLK, Q => 
                           n_1081, QN => n210_port);
   NEXT_REGISTERS_reg_3_45_inst : DLH_X1 port map( G => n11911, D => N4100, Q 
                           => NEXT_REGISTERS_3_45_port);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => N1859, CK => CLK, Q => 
                           n_1082, QN => n211_port);
   NEXT_REGISTERS_reg_3_44_inst : DLH_X1 port map( G => n11911, D => N4099, Q 
                           => NEXT_REGISTERS_3_44_port);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => N1858, CK => CLK, Q => 
                           n_1083, QN => n212_port);
   NEXT_REGISTERS_reg_3_43_inst : DLH_X1 port map( G => n11911, D => N4098, Q 
                           => NEXT_REGISTERS_3_43_port);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => N1857, CK => CLK, Q => 
                           n_1084, QN => n213_port);
   NEXT_REGISTERS_reg_3_42_inst : DLH_X1 port map( G => n11911, D => N4097, Q 
                           => NEXT_REGISTERS_3_42_port);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => N1856, CK => CLK, Q => 
                           n_1085, QN => n214_port);
   NEXT_REGISTERS_reg_3_41_inst : DLH_X1 port map( G => n11912, D => N4096, Q 
                           => NEXT_REGISTERS_3_41_port);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => N1855, CK => CLK, Q => 
                           n_1086, QN => n215_port);
   NEXT_REGISTERS_reg_3_40_inst : DLH_X1 port map( G => n11912, D => N4095, Q 
                           => NEXT_REGISTERS_3_40_port);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => N1854, CK => CLK, Q => 
                           n_1087, QN => n216_port);
   NEXT_REGISTERS_reg_3_39_inst : DLH_X1 port map( G => n11912, D => N4094, Q 
                           => NEXT_REGISTERS_3_39_port);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => N1853, CK => CLK, Q => 
                           n_1088, QN => n217_port);
   NEXT_REGISTERS_reg_3_38_inst : DLH_X1 port map( G => n11912, D => N4093, Q 
                           => NEXT_REGISTERS_3_38_port);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => N1852, CK => CLK, Q => 
                           n_1089, QN => n218_port);
   NEXT_REGISTERS_reg_3_37_inst : DLH_X1 port map( G => n11912, D => N4092, Q 
                           => NEXT_REGISTERS_3_37_port);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => N1851, CK => CLK, Q => 
                           n_1090, QN => n219_port);
   NEXT_REGISTERS_reg_3_36_inst : DLH_X1 port map( G => n11912, D => N4091, Q 
                           => NEXT_REGISTERS_3_36_port);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => N1850, CK => CLK, Q => 
                           n_1091, QN => n220_port);
   NEXT_REGISTERS_reg_3_35_inst : DLH_X1 port map( G => n11912, D => N4090, Q 
                           => NEXT_REGISTERS_3_35_port);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => N1849, CK => CLK, Q => 
                           n_1092, QN => n221_port);
   NEXT_REGISTERS_reg_3_34_inst : DLH_X1 port map( G => n11912, D => N4089, Q 
                           => NEXT_REGISTERS_3_34_port);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => N1848, CK => CLK, Q => 
                           n_1093, QN => n222_port);
   NEXT_REGISTERS_reg_3_33_inst : DLH_X1 port map( G => n11912, D => N4088, Q 
                           => NEXT_REGISTERS_3_33_port);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => N1847, CK => CLK, Q => 
                           n_1094, QN => n223_port);
   NEXT_REGISTERS_reg_3_32_inst : DLH_X1 port map( G => n11912, D => N4087, Q 
                           => NEXT_REGISTERS_3_32_port);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => N1846, CK => CLK, Q => 
                           n_1095, QN => n224_port);
   NEXT_REGISTERS_reg_3_31_inst : DLH_X1 port map( G => n11912, D => N4086, Q 
                           => NEXT_REGISTERS_3_31_port);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => N1845, CK => CLK, Q => 
                           n_1096, QN => n225_port);
   NEXT_REGISTERS_reg_3_30_inst : DLH_X1 port map( G => n11913, D => N4085, Q 
                           => NEXT_REGISTERS_3_30_port);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => N1844, CK => CLK, Q => 
                           n_1097, QN => n226_port);
   NEXT_REGISTERS_reg_3_29_inst : DLH_X1 port map( G => n11913, D => N4084, Q 
                           => NEXT_REGISTERS_3_29_port);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => N1843, CK => CLK, Q => 
                           n_1098, QN => n227_port);
   NEXT_REGISTERS_reg_3_28_inst : DLH_X1 port map( G => n11913, D => N4083, Q 
                           => NEXT_REGISTERS_3_28_port);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => N1842, CK => CLK, Q => 
                           n_1099, QN => n228_port);
   NEXT_REGISTERS_reg_3_27_inst : DLH_X1 port map( G => n11913, D => N4082, Q 
                           => NEXT_REGISTERS_3_27_port);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => N1841, CK => CLK, Q => 
                           n_1100, QN => n229_port);
   NEXT_REGISTERS_reg_3_26_inst : DLH_X1 port map( G => n11913, D => N4081, Q 
                           => NEXT_REGISTERS_3_26_port);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => N1840, CK => CLK, Q => 
                           n_1101, QN => n230_port);
   NEXT_REGISTERS_reg_3_25_inst : DLH_X1 port map( G => n11913, D => N4080, Q 
                           => NEXT_REGISTERS_3_25_port);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => N1839, CK => CLK, Q => 
                           n_1102, QN => n231_port);
   NEXT_REGISTERS_reg_3_24_inst : DLH_X1 port map( G => n11913, D => N4079, Q 
                           => NEXT_REGISTERS_3_24_port);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => N1838, CK => CLK, Q => 
                           n_1103, QN => n232_port);
   NEXT_REGISTERS_reg_3_23_inst : DLH_X1 port map( G => n11913, D => N4078, Q 
                           => NEXT_REGISTERS_3_23_port);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => N1837, CK => CLK, Q => 
                           n_1104, QN => n233_port);
   NEXT_REGISTERS_reg_3_22_inst : DLH_X1 port map( G => n11913, D => N4077, Q 
                           => NEXT_REGISTERS_3_22_port);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => N1836, CK => CLK, Q => 
                           n_1105, QN => n234_port);
   NEXT_REGISTERS_reg_3_21_inst : DLH_X1 port map( G => n11913, D => N4076, Q 
                           => NEXT_REGISTERS_3_21_port);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => N1835, CK => CLK, Q => 
                           n_1106, QN => n235_port);
   NEXT_REGISTERS_reg_3_20_inst : DLH_X1 port map( G => n11913, D => N4075, Q 
                           => NEXT_REGISTERS_3_20_port);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => N1834, CK => CLK, Q => 
                           n_1107, QN => n236_port);
   NEXT_REGISTERS_reg_3_19_inst : DLH_X1 port map( G => n11914, D => N4074, Q 
                           => NEXT_REGISTERS_3_19_port);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => N1833, CK => CLK, Q => 
                           n_1108, QN => n237_port);
   NEXT_REGISTERS_reg_3_18_inst : DLH_X1 port map( G => n11914, D => N4073, Q 
                           => NEXT_REGISTERS_3_18_port);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => N1832, CK => CLK, Q => 
                           n_1109, QN => n238_port);
   NEXT_REGISTERS_reg_3_17_inst : DLH_X1 port map( G => n11914, D => N4072, Q 
                           => NEXT_REGISTERS_3_17_port);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => N1831, CK => CLK, Q => 
                           n_1110, QN => n239_port);
   NEXT_REGISTERS_reg_3_16_inst : DLH_X1 port map( G => n11914, D => N4071, Q 
                           => NEXT_REGISTERS_3_16_port);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => N1830, CK => CLK, Q => 
                           n_1111, QN => n240_port);
   NEXT_REGISTERS_reg_3_15_inst : DLH_X1 port map( G => n11914, D => N4070, Q 
                           => NEXT_REGISTERS_3_15_port);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => N1829, CK => CLK, Q => 
                           n_1112, QN => n241_port);
   NEXT_REGISTERS_reg_3_14_inst : DLH_X1 port map( G => n11914, D => N4069, Q 
                           => NEXT_REGISTERS_3_14_port);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => N1828, CK => CLK, Q => 
                           n_1113, QN => n242_port);
   NEXT_REGISTERS_reg_3_13_inst : DLH_X1 port map( G => n11914, D => N4068, Q 
                           => NEXT_REGISTERS_3_13_port);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => N1827, CK => CLK, Q => 
                           n_1114, QN => n243_port);
   NEXT_REGISTERS_reg_3_12_inst : DLH_X1 port map( G => n11914, D => N4067, Q 
                           => NEXT_REGISTERS_3_12_port);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => N1826, CK => CLK, Q => 
                           n_1115, QN => n244_port);
   NEXT_REGISTERS_reg_3_11_inst : DLH_X1 port map( G => n11914, D => N4066, Q 
                           => NEXT_REGISTERS_3_11_port);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => N1825, CK => CLK, Q => 
                           n_1116, QN => n245_port);
   NEXT_REGISTERS_reg_3_10_inst : DLH_X1 port map( G => n11914, D => N4065, Q 
                           => NEXT_REGISTERS_3_10_port);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => N1824, CK => CLK, Q => 
                           n_1117, QN => n246_port);
   NEXT_REGISTERS_reg_3_9_inst : DLH_X1 port map( G => n11914, D => N4064, Q =>
                           NEXT_REGISTERS_3_9_port);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => N1823, CK => CLK, Q => n_1118
                           , QN => n247_port);
   NEXT_REGISTERS_reg_3_8_inst : DLH_X1 port map( G => n11915, D => N4063, Q =>
                           NEXT_REGISTERS_3_8_port);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => N1822, CK => CLK, Q => n_1119
                           , QN => n248_port);
   NEXT_REGISTERS_reg_3_7_inst : DLH_X1 port map( G => n11915, D => N4062, Q =>
                           NEXT_REGISTERS_3_7_port);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => N1821, CK => CLK, Q => n_1120
                           , QN => n249_port);
   NEXT_REGISTERS_reg_3_6_inst : DLH_X1 port map( G => n11915, D => N4061, Q =>
                           NEXT_REGISTERS_3_6_port);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => N1820, CK => CLK, Q => n_1121
                           , QN => n250_port);
   NEXT_REGISTERS_reg_3_5_inst : DLH_X1 port map( G => n11915, D => N4060, Q =>
                           NEXT_REGISTERS_3_5_port);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => N1819, CK => CLK, Q => n_1122
                           , QN => n251_port);
   NEXT_REGISTERS_reg_3_4_inst : DLH_X1 port map( G => n11915, D => N4059, Q =>
                           NEXT_REGISTERS_3_4_port);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => N1818, CK => CLK, Q => n_1123
                           , QN => n252_port);
   NEXT_REGISTERS_reg_3_3_inst : DLH_X1 port map( G => n11915, D => N4058, Q =>
                           NEXT_REGISTERS_3_3_port);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => N1817, CK => CLK, Q => n_1124
                           , QN => n253_port);
   NEXT_REGISTERS_reg_3_2_inst : DLH_X1 port map( G => n11915, D => N4057, Q =>
                           NEXT_REGISTERS_3_2_port);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => N1816, CK => CLK, Q => n_1125
                           , QN => n254_port);
   NEXT_REGISTERS_reg_3_1_inst : DLH_X1 port map( G => n11915, D => N4056, Q =>
                           NEXT_REGISTERS_3_1_port);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => N1815, CK => CLK, Q => n_1126
                           , QN => n255_port);
   NEXT_REGISTERS_reg_3_0_inst : DLH_X1 port map( G => n11915, D => N4055, Q =>
                           NEXT_REGISTERS_3_0_port);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => N1814, CK => CLK, Q => n_1127
                           , QN => n256_port);
   NEXT_REGISTERS_reg_4_63_inst : DLH_X1 port map( G => n11919, D => N4053, Q 
                           => NEXT_REGISTERS_4_63_port);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => N1813, CK => CLK, Q => 
                           n_1128, QN => n257_port);
   NEXT_REGISTERS_reg_4_62_inst : DLH_X1 port map( G => n11919, D => N4052, Q 
                           => NEXT_REGISTERS_4_62_port);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => N1812, CK => CLK, Q => 
                           n_1129, QN => n258_port);
   NEXT_REGISTERS_reg_4_61_inst : DLH_X1 port map( G => n11919, D => N4051, Q 
                           => NEXT_REGISTERS_4_61_port);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => N1811, CK => CLK, Q => 
                           n_1130, QN => n259_port);
   NEXT_REGISTERS_reg_4_60_inst : DLH_X1 port map( G => n11919, D => N4050, Q 
                           => NEXT_REGISTERS_4_60_port);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => N1810, CK => CLK, Q => 
                           n_1131, QN => n260_port);
   NEXT_REGISTERS_reg_4_59_inst : DLH_X1 port map( G => n11919, D => N4049, Q 
                           => NEXT_REGISTERS_4_59_port);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => N1809, CK => CLK, Q => 
                           n_1132, QN => n261_port);
   NEXT_REGISTERS_reg_4_58_inst : DLH_X1 port map( G => n11919, D => N4048, Q 
                           => NEXT_REGISTERS_4_58_port);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => N1808, CK => CLK, Q => 
                           n_1133, QN => n262_port);
   NEXT_REGISTERS_reg_4_57_inst : DLH_X1 port map( G => n11919, D => N4047, Q 
                           => NEXT_REGISTERS_4_57_port);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => N1807, CK => CLK, Q => 
                           n_1134, QN => n263_port);
   NEXT_REGISTERS_reg_4_56_inst : DLH_X1 port map( G => n11919, D => N4046, Q 
                           => NEXT_REGISTERS_4_56_port);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => N1806, CK => CLK, Q => 
                           n_1135, QN => n264_port);
   NEXT_REGISTERS_reg_4_55_inst : DLH_X1 port map( G => n11919, D => N4045, Q 
                           => NEXT_REGISTERS_4_55_port);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => N1805, CK => CLK, Q => 
                           n_1136, QN => n265_port);
   NEXT_REGISTERS_reg_4_54_inst : DLH_X1 port map( G => n11919, D => N4044, Q 
                           => NEXT_REGISTERS_4_54_port);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => N1804, CK => CLK, Q => 
                           n_1137, QN => n266_port);
   NEXT_REGISTERS_reg_4_53_inst : DLH_X1 port map( G => n11919, D => N4043, Q 
                           => NEXT_REGISTERS_4_53_port);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => N1803, CK => CLK, Q => 
                           n_1138, QN => n267_port);
   NEXT_REGISTERS_reg_4_52_inst : DLH_X1 port map( G => n11920, D => N4042, Q 
                           => NEXT_REGISTERS_4_52_port);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => N1802, CK => CLK, Q => 
                           n_1139, QN => n268_port);
   NEXT_REGISTERS_reg_4_51_inst : DLH_X1 port map( G => n11920, D => N4041, Q 
                           => NEXT_REGISTERS_4_51_port);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => N1801, CK => CLK, Q => 
                           n_1140, QN => n269_port);
   NEXT_REGISTERS_reg_4_50_inst : DLH_X1 port map( G => n11920, D => N4040, Q 
                           => NEXT_REGISTERS_4_50_port);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => N1800, CK => CLK, Q => 
                           n_1141, QN => n270_port);
   NEXT_REGISTERS_reg_4_49_inst : DLH_X1 port map( G => n11920, D => N4039, Q 
                           => NEXT_REGISTERS_4_49_port);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => N1799, CK => CLK, Q => 
                           n_1142, QN => n271_port);
   NEXT_REGISTERS_reg_4_48_inst : DLH_X1 port map( G => n11920, D => N4038, Q 
                           => NEXT_REGISTERS_4_48_port);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => N1798, CK => CLK, Q => 
                           n_1143, QN => n272_port);
   NEXT_REGISTERS_reg_4_47_inst : DLH_X1 port map( G => n11920, D => N4037, Q 
                           => NEXT_REGISTERS_4_47_port);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => N1797, CK => CLK, Q => 
                           n_1144, QN => n273_port);
   NEXT_REGISTERS_reg_4_46_inst : DLH_X1 port map( G => n11920, D => N4036, Q 
                           => NEXT_REGISTERS_4_46_port);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => N1796, CK => CLK, Q => 
                           n_1145, QN => n274_port);
   NEXT_REGISTERS_reg_4_45_inst : DLH_X1 port map( G => n11920, D => N4035, Q 
                           => NEXT_REGISTERS_4_45_port);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => N1795, CK => CLK, Q => 
                           n_1146, QN => n275_port);
   NEXT_REGISTERS_reg_4_44_inst : DLH_X1 port map( G => n11920, D => N4034, Q 
                           => NEXT_REGISTERS_4_44_port);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => N1794, CK => CLK, Q => 
                           n_1147, QN => n276_port);
   NEXT_REGISTERS_reg_4_43_inst : DLH_X1 port map( G => n11920, D => N4033, Q 
                           => NEXT_REGISTERS_4_43_port);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => N1793, CK => CLK, Q => 
                           n_1148, QN => n277_port);
   NEXT_REGISTERS_reg_4_42_inst : DLH_X1 port map( G => n11920, D => N4032, Q 
                           => NEXT_REGISTERS_4_42_port);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => N1792, CK => CLK, Q => 
                           n_1149, QN => n278_port);
   NEXT_REGISTERS_reg_4_41_inst : DLH_X1 port map( G => n11921, D => N4031, Q 
                           => NEXT_REGISTERS_4_41_port);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => N1791, CK => CLK, Q => 
                           n_1150, QN => n279_port);
   NEXT_REGISTERS_reg_4_40_inst : DLH_X1 port map( G => n11921, D => N4030, Q 
                           => NEXT_REGISTERS_4_40_port);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => N1790, CK => CLK, Q => 
                           n_1151, QN => n280_port);
   NEXT_REGISTERS_reg_4_39_inst : DLH_X1 port map( G => n11921, D => N4029, Q 
                           => NEXT_REGISTERS_4_39_port);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => N1789, CK => CLK, Q => 
                           n_1152, QN => n281_port);
   NEXT_REGISTERS_reg_4_38_inst : DLH_X1 port map( G => n11921, D => N4028, Q 
                           => NEXT_REGISTERS_4_38_port);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => N1788, CK => CLK, Q => 
                           n_1153, QN => n282_port);
   NEXT_REGISTERS_reg_4_37_inst : DLH_X1 port map( G => n11921, D => N4027, Q 
                           => NEXT_REGISTERS_4_37_port);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => N1787, CK => CLK, Q => 
                           n_1154, QN => n283_port);
   NEXT_REGISTERS_reg_4_36_inst : DLH_X1 port map( G => n11921, D => N4026, Q 
                           => NEXT_REGISTERS_4_36_port);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => N1786, CK => CLK, Q => 
                           n_1155, QN => n284_port);
   NEXT_REGISTERS_reg_4_35_inst : DLH_X1 port map( G => n11921, D => N4025, Q 
                           => NEXT_REGISTERS_4_35_port);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => N1785, CK => CLK, Q => 
                           n_1156, QN => n285_port);
   NEXT_REGISTERS_reg_4_34_inst : DLH_X1 port map( G => n11921, D => N4024, Q 
                           => NEXT_REGISTERS_4_34_port);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => N1784, CK => CLK, Q => 
                           n_1157, QN => n286_port);
   NEXT_REGISTERS_reg_4_33_inst : DLH_X1 port map( G => n11921, D => N4023, Q 
                           => NEXT_REGISTERS_4_33_port);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => N1783, CK => CLK, Q => 
                           n_1158, QN => n287_port);
   NEXT_REGISTERS_reg_4_32_inst : DLH_X1 port map( G => n11921, D => N4022, Q 
                           => NEXT_REGISTERS_4_32_port);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => N1782, CK => CLK, Q => 
                           n_1159, QN => n288_port);
   NEXT_REGISTERS_reg_4_31_inst : DLH_X1 port map( G => n11921, D => N4021, Q 
                           => NEXT_REGISTERS_4_31_port);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => N1781, CK => CLK, Q => 
                           n_1160, QN => n289_port);
   NEXT_REGISTERS_reg_4_30_inst : DLH_X1 port map( G => n11922, D => N4020, Q 
                           => NEXT_REGISTERS_4_30_port);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => N1780, CK => CLK, Q => 
                           n_1161, QN => n290_port);
   NEXT_REGISTERS_reg_4_29_inst : DLH_X1 port map( G => n11922, D => N4019, Q 
                           => NEXT_REGISTERS_4_29_port);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => N1779, CK => CLK, Q => 
                           n_1162, QN => n291_port);
   NEXT_REGISTERS_reg_4_28_inst : DLH_X1 port map( G => n11922, D => N4018, Q 
                           => NEXT_REGISTERS_4_28_port);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => N1778, CK => CLK, Q => 
                           n_1163, QN => n292_port);
   NEXT_REGISTERS_reg_4_27_inst : DLH_X1 port map( G => n11922, D => N4017, Q 
                           => NEXT_REGISTERS_4_27_port);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => N1777, CK => CLK, Q => 
                           n_1164, QN => n293_port);
   NEXT_REGISTERS_reg_4_26_inst : DLH_X1 port map( G => n11922, D => N4016, Q 
                           => NEXT_REGISTERS_4_26_port);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => N1776, CK => CLK, Q => 
                           n_1165, QN => n294_port);
   NEXT_REGISTERS_reg_4_25_inst : DLH_X1 port map( G => n11922, D => N4015, Q 
                           => NEXT_REGISTERS_4_25_port);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => N1775, CK => CLK, Q => 
                           n_1166, QN => n295_port);
   NEXT_REGISTERS_reg_4_24_inst : DLH_X1 port map( G => n11922, D => N4014, Q 
                           => NEXT_REGISTERS_4_24_port);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => N1774, CK => CLK, Q => 
                           n_1167, QN => n296_port);
   NEXT_REGISTERS_reg_4_23_inst : DLH_X1 port map( G => n11922, D => N4013, Q 
                           => NEXT_REGISTERS_4_23_port);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => N1773, CK => CLK, Q => 
                           n_1168, QN => n297_port);
   NEXT_REGISTERS_reg_4_22_inst : DLH_X1 port map( G => n11922, D => N4012, Q 
                           => NEXT_REGISTERS_4_22_port);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => N1772, CK => CLK, Q => 
                           n_1169, QN => n298_port);
   NEXT_REGISTERS_reg_4_21_inst : DLH_X1 port map( G => n11922, D => N4011, Q 
                           => NEXT_REGISTERS_4_21_port);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => N1771, CK => CLK, Q => 
                           n_1170, QN => n299_port);
   NEXT_REGISTERS_reg_4_20_inst : DLH_X1 port map( G => n11922, D => N4010, Q 
                           => NEXT_REGISTERS_4_20_port);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => N1770, CK => CLK, Q => 
                           n_1171, QN => n300_port);
   NEXT_REGISTERS_reg_4_19_inst : DLH_X1 port map( G => n11923, D => N4009, Q 
                           => NEXT_REGISTERS_4_19_port);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => N1769, CK => CLK, Q => 
                           n_1172, QN => n301_port);
   NEXT_REGISTERS_reg_4_18_inst : DLH_X1 port map( G => n11923, D => N4008, Q 
                           => NEXT_REGISTERS_4_18_port);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => N1768, CK => CLK, Q => 
                           n_1173, QN => n302_port);
   NEXT_REGISTERS_reg_4_17_inst : DLH_X1 port map( G => n11923, D => N4007, Q 
                           => NEXT_REGISTERS_4_17_port);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => N1767, CK => CLK, Q => 
                           n_1174, QN => n303_port);
   NEXT_REGISTERS_reg_4_16_inst : DLH_X1 port map( G => n11923, D => N4006, Q 
                           => NEXT_REGISTERS_4_16_port);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => N1766, CK => CLK, Q => 
                           n_1175, QN => n304_port);
   NEXT_REGISTERS_reg_4_15_inst : DLH_X1 port map( G => n11923, D => N4005, Q 
                           => NEXT_REGISTERS_4_15_port);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => N1765, CK => CLK, Q => 
                           n_1176, QN => n305_port);
   NEXT_REGISTERS_reg_4_14_inst : DLH_X1 port map( G => n11923, D => N4004, Q 
                           => NEXT_REGISTERS_4_14_port);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => N1764, CK => CLK, Q => 
                           n_1177, QN => n306_port);
   NEXT_REGISTERS_reg_4_13_inst : DLH_X1 port map( G => n11923, D => N4003, Q 
                           => NEXT_REGISTERS_4_13_port);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => N1763, CK => CLK, Q => 
                           n_1178, QN => n307_port);
   NEXT_REGISTERS_reg_4_12_inst : DLH_X1 port map( G => n11923, D => N4002, Q 
                           => NEXT_REGISTERS_4_12_port);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => N1762, CK => CLK, Q => 
                           n_1179, QN => n308_port);
   NEXT_REGISTERS_reg_4_11_inst : DLH_X1 port map( G => n11923, D => N4001, Q 
                           => NEXT_REGISTERS_4_11_port);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => N1761, CK => CLK, Q => 
                           n_1180, QN => n309_port);
   NEXT_REGISTERS_reg_4_10_inst : DLH_X1 port map( G => n11923, D => N4000, Q 
                           => NEXT_REGISTERS_4_10_port);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => N1760, CK => CLK, Q => 
                           n_1181, QN => n310_port);
   NEXT_REGISTERS_reg_4_9_inst : DLH_X1 port map( G => n11923, D => N3999, Q =>
                           NEXT_REGISTERS_4_9_port);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => N1759, CK => CLK, Q => n_1182
                           , QN => n311_port);
   NEXT_REGISTERS_reg_4_8_inst : DLH_X1 port map( G => n11924, D => N3998, Q =>
                           NEXT_REGISTERS_4_8_port);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => N1758, CK => CLK, Q => n_1183
                           , QN => n312_port);
   NEXT_REGISTERS_reg_4_7_inst : DLH_X1 port map( G => n11924, D => N3997, Q =>
                           NEXT_REGISTERS_4_7_port);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => N1757, CK => CLK, Q => n_1184
                           , QN => n313_port);
   NEXT_REGISTERS_reg_4_6_inst : DLH_X1 port map( G => n11924, D => N3996, Q =>
                           NEXT_REGISTERS_4_6_port);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => N1756, CK => CLK, Q => n_1185
                           , QN => n314_port);
   NEXT_REGISTERS_reg_4_5_inst : DLH_X1 port map( G => n11924, D => N3995, Q =>
                           NEXT_REGISTERS_4_5_port);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => N1755, CK => CLK, Q => n_1186
                           , QN => n315_port);
   NEXT_REGISTERS_reg_4_4_inst : DLH_X1 port map( G => n11924, D => N3994, Q =>
                           NEXT_REGISTERS_4_4_port);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => N1754, CK => CLK, Q => n_1187
                           , QN => n316_port);
   NEXT_REGISTERS_reg_4_3_inst : DLH_X1 port map( G => n11924, D => N3993, Q =>
                           NEXT_REGISTERS_4_3_port);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => N1753, CK => CLK, Q => n_1188
                           , QN => n317_port);
   NEXT_REGISTERS_reg_4_2_inst : DLH_X1 port map( G => n11924, D => N3992, Q =>
                           NEXT_REGISTERS_4_2_port);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => N1752, CK => CLK, Q => n_1189
                           , QN => n318_port);
   NEXT_REGISTERS_reg_4_1_inst : DLH_X1 port map( G => n11924, D => N3991, Q =>
                           NEXT_REGISTERS_4_1_port);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => N1751, CK => CLK, Q => n_1190
                           , QN => n319_port);
   NEXT_REGISTERS_reg_4_0_inst : DLH_X1 port map( G => n11924, D => N3990, Q =>
                           NEXT_REGISTERS_4_0_port);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => N1750, CK => CLK, Q => n_1191
                           , QN => n320_port);
   NEXT_REGISTERS_reg_5_63_inst : DLH_X1 port map( G => n11928, D => N3988, Q 
                           => NEXT_REGISTERS_5_63_port);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => N1749, CK => CLK, Q => n9965
                           , QN => n321_port);
   NEXT_REGISTERS_reg_5_62_inst : DLH_X1 port map( G => n11928, D => N3987, Q 
                           => NEXT_REGISTERS_5_62_port);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => N1748, CK => CLK, Q => n9963
                           , QN => n322_port);
   NEXT_REGISTERS_reg_5_61_inst : DLH_X1 port map( G => n11928, D => N3986, Q 
                           => NEXT_REGISTERS_5_61_port);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => N1747, CK => CLK, Q => n9961
                           , QN => n323_port);
   NEXT_REGISTERS_reg_5_60_inst : DLH_X1 port map( G => n11928, D => N3985, Q 
                           => NEXT_REGISTERS_5_60_port);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => N1746, CK => CLK, Q => n9959
                           , QN => n324_port);
   NEXT_REGISTERS_reg_5_59_inst : DLH_X1 port map( G => n11928, D => N3984, Q 
                           => NEXT_REGISTERS_5_59_port);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => N1745, CK => CLK, Q => n9957
                           , QN => n325_port);
   NEXT_REGISTERS_reg_5_58_inst : DLH_X1 port map( G => n11928, D => N3983, Q 
                           => NEXT_REGISTERS_5_58_port);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => N1744, CK => CLK, Q => n9955
                           , QN => n326_port);
   NEXT_REGISTERS_reg_5_57_inst : DLH_X1 port map( G => n11928, D => N3982, Q 
                           => NEXT_REGISTERS_5_57_port);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => N1743, CK => CLK, Q => n9953
                           , QN => n327_port);
   NEXT_REGISTERS_reg_5_56_inst : DLH_X1 port map( G => n11928, D => N3981, Q 
                           => NEXT_REGISTERS_5_56_port);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => N1742, CK => CLK, Q => n9951
                           , QN => n328_port);
   NEXT_REGISTERS_reg_5_55_inst : DLH_X1 port map( G => n11928, D => N3980, Q 
                           => NEXT_REGISTERS_5_55_port);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => N1741, CK => CLK, Q => n9949
                           , QN => n329_port);
   NEXT_REGISTERS_reg_5_54_inst : DLH_X1 port map( G => n11928, D => N3979, Q 
                           => NEXT_REGISTERS_5_54_port);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => N1740, CK => CLK, Q => n9947
                           , QN => n330_port);
   NEXT_REGISTERS_reg_5_53_inst : DLH_X1 port map( G => n11928, D => N3978, Q 
                           => NEXT_REGISTERS_5_53_port);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => N1739, CK => CLK, Q => n9945
                           , QN => n331_port);
   NEXT_REGISTERS_reg_5_52_inst : DLH_X1 port map( G => n11929, D => N3977, Q 
                           => NEXT_REGISTERS_5_52_port);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => N1738, CK => CLK, Q => n9943
                           , QN => n332_port);
   NEXT_REGISTERS_reg_5_51_inst : DLH_X1 port map( G => n11929, D => N3976, Q 
                           => NEXT_REGISTERS_5_51_port);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => N1737, CK => CLK, Q => n9941
                           , QN => n333_port);
   NEXT_REGISTERS_reg_5_50_inst : DLH_X1 port map( G => n11929, D => N3975, Q 
                           => NEXT_REGISTERS_5_50_port);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => N1736, CK => CLK, Q => n9939
                           , QN => n334_port);
   NEXT_REGISTERS_reg_5_49_inst : DLH_X1 port map( G => n11929, D => N3974, Q 
                           => NEXT_REGISTERS_5_49_port);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => N1735, CK => CLK, Q => n9937
                           , QN => n335_port);
   NEXT_REGISTERS_reg_5_48_inst : DLH_X1 port map( G => n11929, D => N3973, Q 
                           => NEXT_REGISTERS_5_48_port);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => N1734, CK => CLK, Q => n9935
                           , QN => n336_port);
   NEXT_REGISTERS_reg_5_47_inst : DLH_X1 port map( G => n11929, D => N3972, Q 
                           => NEXT_REGISTERS_5_47_port);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => N1733, CK => CLK, Q => n9933
                           , QN => n337_port);
   NEXT_REGISTERS_reg_5_46_inst : DLH_X1 port map( G => n11929, D => N3971, Q 
                           => NEXT_REGISTERS_5_46_port);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => N1732, CK => CLK, Q => n9931
                           , QN => n338_port);
   NEXT_REGISTERS_reg_5_45_inst : DLH_X1 port map( G => n11929, D => N3970, Q 
                           => NEXT_REGISTERS_5_45_port);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => N1731, CK => CLK, Q => n9929
                           , QN => n339_port);
   NEXT_REGISTERS_reg_5_44_inst : DLH_X1 port map( G => n11929, D => N3969, Q 
                           => NEXT_REGISTERS_5_44_port);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => N1730, CK => CLK, Q => n9927
                           , QN => n340_port);
   NEXT_REGISTERS_reg_5_43_inst : DLH_X1 port map( G => n11929, D => N3968, Q 
                           => NEXT_REGISTERS_5_43_port);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => N1729, CK => CLK, Q => n9925
                           , QN => n341_port);
   NEXT_REGISTERS_reg_5_42_inst : DLH_X1 port map( G => n11929, D => N3967, Q 
                           => NEXT_REGISTERS_5_42_port);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => N1728, CK => CLK, Q => n9923
                           , QN => n342_port);
   NEXT_REGISTERS_reg_5_41_inst : DLH_X1 port map( G => n11930, D => N3966, Q 
                           => NEXT_REGISTERS_5_41_port);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => N1727, CK => CLK, Q => n9921
                           , QN => n343_port);
   NEXT_REGISTERS_reg_5_40_inst : DLH_X1 port map( G => n11930, D => N3965, Q 
                           => NEXT_REGISTERS_5_40_port);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => N1726, CK => CLK, Q => n9919
                           , QN => n344_port);
   NEXT_REGISTERS_reg_5_39_inst : DLH_X1 port map( G => n11930, D => N3964, Q 
                           => NEXT_REGISTERS_5_39_port);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => N1725, CK => CLK, Q => n9917
                           , QN => n345_port);
   NEXT_REGISTERS_reg_5_38_inst : DLH_X1 port map( G => n11930, D => N3963, Q 
                           => NEXT_REGISTERS_5_38_port);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => N1724, CK => CLK, Q => n9915
                           , QN => n346_port);
   NEXT_REGISTERS_reg_5_37_inst : DLH_X1 port map( G => n11930, D => N3962, Q 
                           => NEXT_REGISTERS_5_37_port);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => N1723, CK => CLK, Q => n9913
                           , QN => n347_port);
   NEXT_REGISTERS_reg_5_36_inst : DLH_X1 port map( G => n11930, D => N3961, Q 
                           => NEXT_REGISTERS_5_36_port);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => N1722, CK => CLK, Q => n9911
                           , QN => n348_port);
   NEXT_REGISTERS_reg_5_35_inst : DLH_X1 port map( G => n11930, D => N3960, Q 
                           => NEXT_REGISTERS_5_35_port);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => N1721, CK => CLK, Q => n9909
                           , QN => n349_port);
   NEXT_REGISTERS_reg_5_34_inst : DLH_X1 port map( G => n11930, D => N3959, Q 
                           => NEXT_REGISTERS_5_34_port);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => N1720, CK => CLK, Q => n9907
                           , QN => n350_port);
   NEXT_REGISTERS_reg_5_33_inst : DLH_X1 port map( G => n11930, D => N3958, Q 
                           => NEXT_REGISTERS_5_33_port);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => N1719, CK => CLK, Q => n9905
                           , QN => n351_port);
   NEXT_REGISTERS_reg_5_32_inst : DLH_X1 port map( G => n11930, D => N3957, Q 
                           => NEXT_REGISTERS_5_32_port);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => N1718, CK => CLK, Q => n9903
                           , QN => n352_port);
   NEXT_REGISTERS_reg_5_31_inst : DLH_X1 port map( G => n11930, D => N3956, Q 
                           => NEXT_REGISTERS_5_31_port);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => N1717, CK => CLK, Q => n9901
                           , QN => n353_port);
   NEXT_REGISTERS_reg_5_30_inst : DLH_X1 port map( G => n11931, D => N3955, Q 
                           => NEXT_REGISTERS_5_30_port);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => N1716, CK => CLK, Q => n9899
                           , QN => n354_port);
   NEXT_REGISTERS_reg_5_29_inst : DLH_X1 port map( G => n11931, D => N3954, Q 
                           => NEXT_REGISTERS_5_29_port);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => N1715, CK => CLK, Q => n9897
                           , QN => n355_port);
   NEXT_REGISTERS_reg_5_28_inst : DLH_X1 port map( G => n11931, D => N3953, Q 
                           => NEXT_REGISTERS_5_28_port);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => N1714, CK => CLK, Q => n9895
                           , QN => n356_port);
   NEXT_REGISTERS_reg_5_27_inst : DLH_X1 port map( G => n11931, D => N3952, Q 
                           => NEXT_REGISTERS_5_27_port);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => N1713, CK => CLK, Q => n9893
                           , QN => n357_port);
   NEXT_REGISTERS_reg_5_26_inst : DLH_X1 port map( G => n11931, D => N3951, Q 
                           => NEXT_REGISTERS_5_26_port);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => N1712, CK => CLK, Q => n9891
                           , QN => n358_port);
   NEXT_REGISTERS_reg_5_25_inst : DLH_X1 port map( G => n11931, D => N3950, Q 
                           => NEXT_REGISTERS_5_25_port);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => N1711, CK => CLK, Q => n9889
                           , QN => n359_port);
   NEXT_REGISTERS_reg_5_24_inst : DLH_X1 port map( G => n11931, D => N3949, Q 
                           => NEXT_REGISTERS_5_24_port);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => N1710, CK => CLK, Q => n9887
                           , QN => n360_port);
   NEXT_REGISTERS_reg_5_23_inst : DLH_X1 port map( G => n11931, D => N3948, Q 
                           => NEXT_REGISTERS_5_23_port);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => N1709, CK => CLK, Q => n9885
                           , QN => n361_port);
   NEXT_REGISTERS_reg_5_22_inst : DLH_X1 port map( G => n11931, D => N3947, Q 
                           => NEXT_REGISTERS_5_22_port);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => N1708, CK => CLK, Q => n9883
                           , QN => n362_port);
   NEXT_REGISTERS_reg_5_21_inst : DLH_X1 port map( G => n11931, D => N3946, Q 
                           => NEXT_REGISTERS_5_21_port);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => N1707, CK => CLK, Q => n9881
                           , QN => n363_port);
   NEXT_REGISTERS_reg_5_20_inst : DLH_X1 port map( G => n11931, D => N3945, Q 
                           => NEXT_REGISTERS_5_20_port);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => N1706, CK => CLK, Q => n9879
                           , QN => n364_port);
   NEXT_REGISTERS_reg_5_19_inst : DLH_X1 port map( G => n11932, D => N3944, Q 
                           => NEXT_REGISTERS_5_19_port);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => N1705, CK => CLK, Q => n9877
                           , QN => n365_port);
   NEXT_REGISTERS_reg_5_18_inst : DLH_X1 port map( G => n11932, D => N3943, Q 
                           => NEXT_REGISTERS_5_18_port);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => N1704, CK => CLK, Q => n9875
                           , QN => n366_port);
   NEXT_REGISTERS_reg_5_17_inst : DLH_X1 port map( G => n11932, D => N3942, Q 
                           => NEXT_REGISTERS_5_17_port);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => N1703, CK => CLK, Q => n9873
                           , QN => n367_port);
   NEXT_REGISTERS_reg_5_16_inst : DLH_X1 port map( G => n11932, D => N3941, Q 
                           => NEXT_REGISTERS_5_16_port);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => N1702, CK => CLK, Q => n9871
                           , QN => n368_port);
   NEXT_REGISTERS_reg_5_15_inst : DLH_X1 port map( G => n11932, D => N3940, Q 
                           => NEXT_REGISTERS_5_15_port);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => N1701, CK => CLK, Q => n9869
                           , QN => n369_port);
   NEXT_REGISTERS_reg_5_14_inst : DLH_X1 port map( G => n11932, D => N3939, Q 
                           => NEXT_REGISTERS_5_14_port);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => N1700, CK => CLK, Q => n9867
                           , QN => n370_port);
   NEXT_REGISTERS_reg_5_13_inst : DLH_X1 port map( G => n11932, D => N3938, Q 
                           => NEXT_REGISTERS_5_13_port);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => N1699, CK => CLK, Q => n9865
                           , QN => n371_port);
   NEXT_REGISTERS_reg_5_12_inst : DLH_X1 port map( G => n11932, D => N3937, Q 
                           => NEXT_REGISTERS_5_12_port);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => N1698, CK => CLK, Q => n9863
                           , QN => n372_port);
   NEXT_REGISTERS_reg_5_11_inst : DLH_X1 port map( G => n11932, D => N3936, Q 
                           => NEXT_REGISTERS_5_11_port);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => N1697, CK => CLK, Q => n9861
                           , QN => n373_port);
   NEXT_REGISTERS_reg_5_10_inst : DLH_X1 port map( G => n11932, D => N3935, Q 
                           => NEXT_REGISTERS_5_10_port);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => N1696, CK => CLK, Q => n9859
                           , QN => n374_port);
   NEXT_REGISTERS_reg_5_9_inst : DLH_X1 port map( G => n11932, D => N3934, Q =>
                           NEXT_REGISTERS_5_9_port);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => N1695, CK => CLK, Q => n9857,
                           QN => n375_port);
   NEXT_REGISTERS_reg_5_8_inst : DLH_X1 port map( G => n11933, D => N3933, Q =>
                           NEXT_REGISTERS_5_8_port);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => N1694, CK => CLK, Q => n9855,
                           QN => n376_port);
   NEXT_REGISTERS_reg_5_7_inst : DLH_X1 port map( G => n11933, D => N3932, Q =>
                           NEXT_REGISTERS_5_7_port);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => N1693, CK => CLK, Q => n9853,
                           QN => n377_port);
   NEXT_REGISTERS_reg_5_6_inst : DLH_X1 port map( G => n11933, D => N3931, Q =>
                           NEXT_REGISTERS_5_6_port);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => N1692, CK => CLK, Q => n9851,
                           QN => n378_port);
   NEXT_REGISTERS_reg_5_5_inst : DLH_X1 port map( G => n11933, D => N3930, Q =>
                           NEXT_REGISTERS_5_5_port);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => N1691, CK => CLK, Q => n9849,
                           QN => n379_port);
   NEXT_REGISTERS_reg_5_4_inst : DLH_X1 port map( G => n11933, D => N3929, Q =>
                           NEXT_REGISTERS_5_4_port);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => N1690, CK => CLK, Q => n9847,
                           QN => n380_port);
   NEXT_REGISTERS_reg_5_3_inst : DLH_X1 port map( G => n11933, D => N3928, Q =>
                           NEXT_REGISTERS_5_3_port);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => N1689, CK => CLK, Q => n9845,
                           QN => n381_port);
   NEXT_REGISTERS_reg_5_2_inst : DLH_X1 port map( G => n11933, D => N3927, Q =>
                           NEXT_REGISTERS_5_2_port);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => N1688, CK => CLK, Q => n9843,
                           QN => n382_port);
   NEXT_REGISTERS_reg_5_1_inst : DLH_X1 port map( G => n11933, D => N3926, Q =>
                           NEXT_REGISTERS_5_1_port);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => N1687, CK => CLK, Q => n9841,
                           QN => n383_port);
   NEXT_REGISTERS_reg_5_0_inst : DLH_X1 port map( G => n11933, D => N3925, Q =>
                           NEXT_REGISTERS_5_0_port);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => N1686, CK => CLK, Q => n9839,
                           QN => n384_port);
   NEXT_REGISTERS_reg_6_63_inst : DLH_X1 port map( G => n11937, D => N3923, Q 
                           => NEXT_REGISTERS_6_63_port);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => N1685, CK => CLK, Q => 
                           n_1192, QN => n385_port);
   NEXT_REGISTERS_reg_6_62_inst : DLH_X1 port map( G => n11937, D => N3922, Q 
                           => NEXT_REGISTERS_6_62_port);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => N1684, CK => CLK, Q => 
                           n_1193, QN => n386_port);
   NEXT_REGISTERS_reg_6_61_inst : DLH_X1 port map( G => n11937, D => N3921, Q 
                           => NEXT_REGISTERS_6_61_port);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => N1683, CK => CLK, Q => 
                           n_1194, QN => n387_port);
   NEXT_REGISTERS_reg_6_60_inst : DLH_X1 port map( G => n11937, D => N3920, Q 
                           => NEXT_REGISTERS_6_60_port);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => N1682, CK => CLK, Q => 
                           n_1195, QN => n388_port);
   NEXT_REGISTERS_reg_6_59_inst : DLH_X1 port map( G => n11937, D => N3919, Q 
                           => NEXT_REGISTERS_6_59_port);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => N1681, CK => CLK, Q => 
                           n_1196, QN => n389_port);
   NEXT_REGISTERS_reg_6_58_inst : DLH_X1 port map( G => n11937, D => N3918, Q 
                           => NEXT_REGISTERS_6_58_port);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => N1680, CK => CLK, Q => 
                           n_1197, QN => n390_port);
   NEXT_REGISTERS_reg_6_57_inst : DLH_X1 port map( G => n11937, D => N3917, Q 
                           => NEXT_REGISTERS_6_57_port);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => N1679, CK => CLK, Q => 
                           n_1198, QN => n391_port);
   NEXT_REGISTERS_reg_6_56_inst : DLH_X1 port map( G => n11937, D => N3916, Q 
                           => NEXT_REGISTERS_6_56_port);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => N1678, CK => CLK, Q => 
                           n_1199, QN => n392_port);
   NEXT_REGISTERS_reg_6_55_inst : DLH_X1 port map( G => n11937, D => N3915, Q 
                           => NEXT_REGISTERS_6_55_port);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => N1677, CK => CLK, Q => 
                           n_1200, QN => n393_port);
   NEXT_REGISTERS_reg_6_54_inst : DLH_X1 port map( G => n11937, D => N3914, Q 
                           => NEXT_REGISTERS_6_54_port);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => N1676, CK => CLK, Q => 
                           n_1201, QN => n394_port);
   NEXT_REGISTERS_reg_6_53_inst : DLH_X1 port map( G => n11937, D => N3913, Q 
                           => NEXT_REGISTERS_6_53_port);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => N1675, CK => CLK, Q => 
                           n_1202, QN => n395_port);
   NEXT_REGISTERS_reg_6_52_inst : DLH_X1 port map( G => n11938, D => N3912, Q 
                           => NEXT_REGISTERS_6_52_port);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => N1674, CK => CLK, Q => 
                           n_1203, QN => n396_port);
   NEXT_REGISTERS_reg_6_51_inst : DLH_X1 port map( G => n11938, D => N3911, Q 
                           => NEXT_REGISTERS_6_51_port);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => N1673, CK => CLK, Q => 
                           n_1204, QN => n397_port);
   NEXT_REGISTERS_reg_6_50_inst : DLH_X1 port map( G => n11938, D => N3910, Q 
                           => NEXT_REGISTERS_6_50_port);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => N1672, CK => CLK, Q => 
                           n_1205, QN => n398_port);
   NEXT_REGISTERS_reg_6_49_inst : DLH_X1 port map( G => n11938, D => N3909, Q 
                           => NEXT_REGISTERS_6_49_port);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => N1671, CK => CLK, Q => 
                           n_1206, QN => n399_port);
   NEXT_REGISTERS_reg_6_48_inst : DLH_X1 port map( G => n11938, D => N3908, Q 
                           => NEXT_REGISTERS_6_48_port);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => N1670, CK => CLK, Q => 
                           n_1207, QN => n400_port);
   NEXT_REGISTERS_reg_6_47_inst : DLH_X1 port map( G => n11938, D => N3907, Q 
                           => NEXT_REGISTERS_6_47_port);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => N1669, CK => CLK, Q => 
                           n_1208, QN => n401_port);
   NEXT_REGISTERS_reg_6_46_inst : DLH_X1 port map( G => n11938, D => N3906, Q 
                           => NEXT_REGISTERS_6_46_port);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => N1668, CK => CLK, Q => 
                           n_1209, QN => n402_port);
   NEXT_REGISTERS_reg_6_45_inst : DLH_X1 port map( G => n11938, D => N3905, Q 
                           => NEXT_REGISTERS_6_45_port);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => N1667, CK => CLK, Q => 
                           n_1210, QN => n403_port);
   NEXT_REGISTERS_reg_6_44_inst : DLH_X1 port map( G => n11938, D => N3904, Q 
                           => NEXT_REGISTERS_6_44_port);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => N1666, CK => CLK, Q => 
                           n_1211, QN => n404_port);
   NEXT_REGISTERS_reg_6_43_inst : DLH_X1 port map( G => n11938, D => N3903, Q 
                           => NEXT_REGISTERS_6_43_port);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => N1665, CK => CLK, Q => 
                           n_1212, QN => n405_port);
   NEXT_REGISTERS_reg_6_42_inst : DLH_X1 port map( G => n11938, D => N3902, Q 
                           => NEXT_REGISTERS_6_42_port);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => N1664, CK => CLK, Q => 
                           n_1213, QN => n406_port);
   NEXT_REGISTERS_reg_6_41_inst : DLH_X1 port map( G => n11939, D => N3901, Q 
                           => NEXT_REGISTERS_6_41_port);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => N1663, CK => CLK, Q => 
                           n_1214, QN => n407_port);
   NEXT_REGISTERS_reg_6_40_inst : DLH_X1 port map( G => n11939, D => N3900, Q 
                           => NEXT_REGISTERS_6_40_port);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => N1662, CK => CLK, Q => 
                           n_1215, QN => n408_port);
   NEXT_REGISTERS_reg_6_39_inst : DLH_X1 port map( G => n11939, D => N3899, Q 
                           => NEXT_REGISTERS_6_39_port);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => N1661, CK => CLK, Q => 
                           n_1216, QN => n409_port);
   NEXT_REGISTERS_reg_6_38_inst : DLH_X1 port map( G => n11939, D => N3898, Q 
                           => NEXT_REGISTERS_6_38_port);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => N1660, CK => CLK, Q => 
                           n_1217, QN => n410_port);
   NEXT_REGISTERS_reg_6_37_inst : DLH_X1 port map( G => n11939, D => N3897, Q 
                           => NEXT_REGISTERS_6_37_port);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => N1659, CK => CLK, Q => 
                           n_1218, QN => n411_port);
   NEXT_REGISTERS_reg_6_36_inst : DLH_X1 port map( G => n11939, D => N3896, Q 
                           => NEXT_REGISTERS_6_36_port);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => N1658, CK => CLK, Q => 
                           n_1219, QN => n412_port);
   NEXT_REGISTERS_reg_6_35_inst : DLH_X1 port map( G => n11939, D => N3895, Q 
                           => NEXT_REGISTERS_6_35_port);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => N1657, CK => CLK, Q => 
                           n_1220, QN => n413_port);
   NEXT_REGISTERS_reg_6_34_inst : DLH_X1 port map( G => n11939, D => N3894, Q 
                           => NEXT_REGISTERS_6_34_port);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => N1656, CK => CLK, Q => 
                           n_1221, QN => n414_port);
   NEXT_REGISTERS_reg_6_33_inst : DLH_X1 port map( G => n11939, D => N3893, Q 
                           => NEXT_REGISTERS_6_33_port);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => N1655, CK => CLK, Q => 
                           n_1222, QN => n415_port);
   NEXT_REGISTERS_reg_6_32_inst : DLH_X1 port map( G => n11939, D => N3892, Q 
                           => NEXT_REGISTERS_6_32_port);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => N1654, CK => CLK, Q => 
                           n_1223, QN => n416_port);
   NEXT_REGISTERS_reg_6_31_inst : DLH_X1 port map( G => n11939, D => N3891, Q 
                           => NEXT_REGISTERS_6_31_port);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => N1653, CK => CLK, Q => 
                           n_1224, QN => n417_port);
   NEXT_REGISTERS_reg_6_30_inst : DLH_X1 port map( G => n11940, D => N3890, Q 
                           => NEXT_REGISTERS_6_30_port);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => N1652, CK => CLK, Q => 
                           n_1225, QN => n418_port);
   NEXT_REGISTERS_reg_6_29_inst : DLH_X1 port map( G => n11940, D => N3889, Q 
                           => NEXT_REGISTERS_6_29_port);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => N1651, CK => CLK, Q => 
                           n_1226, QN => n419_port);
   NEXT_REGISTERS_reg_6_28_inst : DLH_X1 port map( G => n11940, D => N3888, Q 
                           => NEXT_REGISTERS_6_28_port);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => N1650, CK => CLK, Q => 
                           n_1227, QN => n420_port);
   NEXT_REGISTERS_reg_6_27_inst : DLH_X1 port map( G => n11940, D => N3887, Q 
                           => NEXT_REGISTERS_6_27_port);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => N1649, CK => CLK, Q => 
                           n_1228, QN => n421_port);
   NEXT_REGISTERS_reg_6_26_inst : DLH_X1 port map( G => n11940, D => N3886, Q 
                           => NEXT_REGISTERS_6_26_port);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => N1648, CK => CLK, Q => 
                           n_1229, QN => n422_port);
   NEXT_REGISTERS_reg_6_25_inst : DLH_X1 port map( G => n11940, D => N3885, Q 
                           => NEXT_REGISTERS_6_25_port);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => N1647, CK => CLK, Q => 
                           n_1230, QN => n423_port);
   NEXT_REGISTERS_reg_6_24_inst : DLH_X1 port map( G => n11940, D => N3884, Q 
                           => NEXT_REGISTERS_6_24_port);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => N1646, CK => CLK, Q => 
                           n_1231, QN => n424_port);
   NEXT_REGISTERS_reg_6_23_inst : DLH_X1 port map( G => n11940, D => N3883, Q 
                           => NEXT_REGISTERS_6_23_port);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => N1645, CK => CLK, Q => 
                           n_1232, QN => n425_port);
   NEXT_REGISTERS_reg_6_22_inst : DLH_X1 port map( G => n11940, D => N3882, Q 
                           => NEXT_REGISTERS_6_22_port);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => N1644, CK => CLK, Q => 
                           n_1233, QN => n426_port);
   NEXT_REGISTERS_reg_6_21_inst : DLH_X1 port map( G => n11940, D => N3881, Q 
                           => NEXT_REGISTERS_6_21_port);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => N1643, CK => CLK, Q => 
                           n_1234, QN => n427_port);
   NEXT_REGISTERS_reg_6_20_inst : DLH_X1 port map( G => n11940, D => N3880, Q 
                           => NEXT_REGISTERS_6_20_port);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => N1642, CK => CLK, Q => 
                           n_1235, QN => n428_port);
   NEXT_REGISTERS_reg_6_19_inst : DLH_X1 port map( G => n11941, D => N3879, Q 
                           => NEXT_REGISTERS_6_19_port);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => N1641, CK => CLK, Q => 
                           n_1236, QN => n429_port);
   NEXT_REGISTERS_reg_6_18_inst : DLH_X1 port map( G => n11941, D => N3878, Q 
                           => NEXT_REGISTERS_6_18_port);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => N1640, CK => CLK, Q => 
                           n_1237, QN => n430_port);
   NEXT_REGISTERS_reg_6_17_inst : DLH_X1 port map( G => n11941, D => N3877, Q 
                           => NEXT_REGISTERS_6_17_port);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => N1639, CK => CLK, Q => 
                           n_1238, QN => n431_port);
   NEXT_REGISTERS_reg_6_16_inst : DLH_X1 port map( G => n11941, D => N3876, Q 
                           => NEXT_REGISTERS_6_16_port);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => N1638, CK => CLK, Q => 
                           n_1239, QN => n432_port);
   NEXT_REGISTERS_reg_6_15_inst : DLH_X1 port map( G => n11941, D => N3875, Q 
                           => NEXT_REGISTERS_6_15_port);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => N1637, CK => CLK, Q => 
                           n_1240, QN => n433_port);
   NEXT_REGISTERS_reg_6_14_inst : DLH_X1 port map( G => n11941, D => N3874, Q 
                           => NEXT_REGISTERS_6_14_port);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => N1636, CK => CLK, Q => 
                           n_1241, QN => n434_port);
   NEXT_REGISTERS_reg_6_13_inst : DLH_X1 port map( G => n11941, D => N3873, Q 
                           => NEXT_REGISTERS_6_13_port);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => N1635, CK => CLK, Q => 
                           n_1242, QN => n435_port);
   NEXT_REGISTERS_reg_6_12_inst : DLH_X1 port map( G => n11941, D => N3872, Q 
                           => NEXT_REGISTERS_6_12_port);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => N1634, CK => CLK, Q => 
                           n_1243, QN => n436_port);
   NEXT_REGISTERS_reg_6_11_inst : DLH_X1 port map( G => n11941, D => N3871, Q 
                           => NEXT_REGISTERS_6_11_port);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => N1633, CK => CLK, Q => 
                           n_1244, QN => n437_port);
   NEXT_REGISTERS_reg_6_10_inst : DLH_X1 port map( G => n11941, D => N3870, Q 
                           => NEXT_REGISTERS_6_10_port);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => N1632, CK => CLK, Q => 
                           n_1245, QN => n438_port);
   NEXT_REGISTERS_reg_6_9_inst : DLH_X1 port map( G => n11941, D => N3869, Q =>
                           NEXT_REGISTERS_6_9_port);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => N1631, CK => CLK, Q => n_1246
                           , QN => n439_port);
   NEXT_REGISTERS_reg_6_8_inst : DLH_X1 port map( G => n11942, D => N3868, Q =>
                           NEXT_REGISTERS_6_8_port);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => N1630, CK => CLK, Q => n_1247
                           , QN => n440_port);
   NEXT_REGISTERS_reg_6_7_inst : DLH_X1 port map( G => n11942, D => N3867, Q =>
                           NEXT_REGISTERS_6_7_port);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => N1629, CK => CLK, Q => n_1248
                           , QN => n441_port);
   NEXT_REGISTERS_reg_6_6_inst : DLH_X1 port map( G => n11942, D => N3866, Q =>
                           NEXT_REGISTERS_6_6_port);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => N1628, CK => CLK, Q => n_1249
                           , QN => n442_port);
   NEXT_REGISTERS_reg_6_5_inst : DLH_X1 port map( G => n11942, D => N3865, Q =>
                           NEXT_REGISTERS_6_5_port);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => N1627, CK => CLK, Q => n_1250
                           , QN => n443_port);
   NEXT_REGISTERS_reg_6_4_inst : DLH_X1 port map( G => n11942, D => N3864, Q =>
                           NEXT_REGISTERS_6_4_port);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => N1626, CK => CLK, Q => n_1251
                           , QN => n444_port);
   NEXT_REGISTERS_reg_6_3_inst : DLH_X1 port map( G => n11942, D => N3863, Q =>
                           NEXT_REGISTERS_6_3_port);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => N1625, CK => CLK, Q => n_1252
                           , QN => n445_port);
   NEXT_REGISTERS_reg_6_2_inst : DLH_X1 port map( G => n11942, D => N3862, Q =>
                           NEXT_REGISTERS_6_2_port);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => N1624, CK => CLK, Q => n_1253
                           , QN => n446_port);
   NEXT_REGISTERS_reg_6_1_inst : DLH_X1 port map( G => n11942, D => N3861, Q =>
                           NEXT_REGISTERS_6_1_port);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => N1623, CK => CLK, Q => n_1254
                           , QN => n447_port);
   NEXT_REGISTERS_reg_6_0_inst : DLH_X1 port map( G => n11942, D => N3860, Q =>
                           NEXT_REGISTERS_6_0_port);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => N1622, CK => CLK, Q => n_1255
                           , QN => n448_port);
   NEXT_REGISTERS_reg_7_63_inst : DLH_X1 port map( G => n11946, D => N3858, Q 
                           => NEXT_REGISTERS_7_63_port);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => N1621, CK => CLK, Q => 
                           n10413, QN => n449_port);
   NEXT_REGISTERS_reg_7_62_inst : DLH_X1 port map( G => n11946, D => N3857, Q 
                           => NEXT_REGISTERS_7_62_port);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => N1620, CK => CLK, Q => 
                           n10411, QN => n450_port);
   NEXT_REGISTERS_reg_7_61_inst : DLH_X1 port map( G => n11946, D => N3856, Q 
                           => NEXT_REGISTERS_7_61_port);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => N1619, CK => CLK, Q => 
                           n10409, QN => n451_port);
   NEXT_REGISTERS_reg_7_60_inst : DLH_X1 port map( G => n11946, D => N3855, Q 
                           => NEXT_REGISTERS_7_60_port);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => N1618, CK => CLK, Q => 
                           n10407, QN => n452_port);
   NEXT_REGISTERS_reg_7_59_inst : DLH_X1 port map( G => n11946, D => N3854, Q 
                           => NEXT_REGISTERS_7_59_port);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => N1617, CK => CLK, Q => 
                           n10405, QN => n453_port);
   NEXT_REGISTERS_reg_7_58_inst : DLH_X1 port map( G => n11946, D => N3853, Q 
                           => NEXT_REGISTERS_7_58_port);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => N1616, CK => CLK, Q => 
                           n10403, QN => n454_port);
   NEXT_REGISTERS_reg_7_57_inst : DLH_X1 port map( G => n11946, D => N3852, Q 
                           => NEXT_REGISTERS_7_57_port);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => N1615, CK => CLK, Q => 
                           n10401, QN => n455_port);
   NEXT_REGISTERS_reg_7_56_inst : DLH_X1 port map( G => n11946, D => N3851, Q 
                           => NEXT_REGISTERS_7_56_port);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => N1614, CK => CLK, Q => 
                           n10399, QN => n456_port);
   NEXT_REGISTERS_reg_7_55_inst : DLH_X1 port map( G => n11946, D => N3850, Q 
                           => NEXT_REGISTERS_7_55_port);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => N1613, CK => CLK, Q => 
                           n10397, QN => n457_port);
   NEXT_REGISTERS_reg_7_54_inst : DLH_X1 port map( G => n11946, D => N3849, Q 
                           => NEXT_REGISTERS_7_54_port);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => N1612, CK => CLK, Q => 
                           n10395, QN => n458_port);
   NEXT_REGISTERS_reg_7_53_inst : DLH_X1 port map( G => n11946, D => N3848, Q 
                           => NEXT_REGISTERS_7_53_port);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => N1611, CK => CLK, Q => 
                           n10393, QN => n459_port);
   NEXT_REGISTERS_reg_7_52_inst : DLH_X1 port map( G => n11947, D => N3847, Q 
                           => NEXT_REGISTERS_7_52_port);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => N1610, CK => CLK, Q => 
                           n10391, QN => n460_port);
   NEXT_REGISTERS_reg_7_51_inst : DLH_X1 port map( G => n11947, D => N3846, Q 
                           => NEXT_REGISTERS_7_51_port);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => N1609, CK => CLK, Q => 
                           n10389, QN => n461_port);
   NEXT_REGISTERS_reg_7_50_inst : DLH_X1 port map( G => n11947, D => N3845, Q 
                           => NEXT_REGISTERS_7_50_port);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => N1608, CK => CLK, Q => 
                           n10387, QN => n462_port);
   NEXT_REGISTERS_reg_7_49_inst : DLH_X1 port map( G => n11947, D => N3844, Q 
                           => NEXT_REGISTERS_7_49_port);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => N1607, CK => CLK, Q => 
                           n10385, QN => n463_port);
   NEXT_REGISTERS_reg_7_48_inst : DLH_X1 port map( G => n11947, D => N3843, Q 
                           => NEXT_REGISTERS_7_48_port);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => N1606, CK => CLK, Q => 
                           n10383, QN => n464_port);
   NEXT_REGISTERS_reg_7_47_inst : DLH_X1 port map( G => n11947, D => N3842, Q 
                           => NEXT_REGISTERS_7_47_port);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => N1605, CK => CLK, Q => 
                           n10381, QN => n465_port);
   NEXT_REGISTERS_reg_7_46_inst : DLH_X1 port map( G => n11947, D => N3841, Q 
                           => NEXT_REGISTERS_7_46_port);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => N1604, CK => CLK, Q => 
                           n10379, QN => n466_port);
   NEXT_REGISTERS_reg_7_45_inst : DLH_X1 port map( G => n11947, D => N3840, Q 
                           => NEXT_REGISTERS_7_45_port);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => N1603, CK => CLK, Q => 
                           n10377, QN => n467_port);
   NEXT_REGISTERS_reg_7_44_inst : DLH_X1 port map( G => n11947, D => N3839, Q 
                           => NEXT_REGISTERS_7_44_port);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => N1602, CK => CLK, Q => 
                           n10375, QN => n468_port);
   NEXT_REGISTERS_reg_7_43_inst : DLH_X1 port map( G => n11947, D => N3838, Q 
                           => NEXT_REGISTERS_7_43_port);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => N1601, CK => CLK, Q => 
                           n10373, QN => n469_port);
   NEXT_REGISTERS_reg_7_42_inst : DLH_X1 port map( G => n11947, D => N3837, Q 
                           => NEXT_REGISTERS_7_42_port);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => N1600, CK => CLK, Q => 
                           n10371, QN => n470_port);
   NEXT_REGISTERS_reg_7_41_inst : DLH_X1 port map( G => n11948, D => N3836, Q 
                           => NEXT_REGISTERS_7_41_port);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => N1599, CK => CLK, Q => 
                           n10369, QN => n471_port);
   NEXT_REGISTERS_reg_7_40_inst : DLH_X1 port map( G => n11948, D => N3835, Q 
                           => NEXT_REGISTERS_7_40_port);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => N1598, CK => CLK, Q => 
                           n10367, QN => n472_port);
   NEXT_REGISTERS_reg_7_39_inst : DLH_X1 port map( G => n11948, D => N3834, Q 
                           => NEXT_REGISTERS_7_39_port);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => N1597, CK => CLK, Q => 
                           n10365, QN => n473_port);
   NEXT_REGISTERS_reg_7_38_inst : DLH_X1 port map( G => n11948, D => N3833, Q 
                           => NEXT_REGISTERS_7_38_port);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => N1596, CK => CLK, Q => 
                           n10363, QN => n474_port);
   NEXT_REGISTERS_reg_7_37_inst : DLH_X1 port map( G => n11948, D => N3832, Q 
                           => NEXT_REGISTERS_7_37_port);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => N1595, CK => CLK, Q => 
                           n10361, QN => n475_port);
   NEXT_REGISTERS_reg_7_36_inst : DLH_X1 port map( G => n11948, D => N3831, Q 
                           => NEXT_REGISTERS_7_36_port);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => N1594, CK => CLK, Q => 
                           n10359, QN => n476_port);
   NEXT_REGISTERS_reg_7_35_inst : DLH_X1 port map( G => n11948, D => N3830, Q 
                           => NEXT_REGISTERS_7_35_port);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => N1593, CK => CLK, Q => 
                           n10357, QN => n477_port);
   NEXT_REGISTERS_reg_7_34_inst : DLH_X1 port map( G => n11948, D => N3829, Q 
                           => NEXT_REGISTERS_7_34_port);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => N1592, CK => CLK, Q => 
                           n10355, QN => n478_port);
   NEXT_REGISTERS_reg_7_33_inst : DLH_X1 port map( G => n11948, D => N3828, Q 
                           => NEXT_REGISTERS_7_33_port);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => N1591, CK => CLK, Q => 
                           n10353, QN => n479_port);
   NEXT_REGISTERS_reg_7_32_inst : DLH_X1 port map( G => n11948, D => N3827, Q 
                           => NEXT_REGISTERS_7_32_port);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => N1590, CK => CLK, Q => 
                           n10351, QN => n480_port);
   NEXT_REGISTERS_reg_7_31_inst : DLH_X1 port map( G => n11948, D => N3826, Q 
                           => NEXT_REGISTERS_7_31_port);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => N1589, CK => CLK, Q => 
                           n10349, QN => n481_port);
   NEXT_REGISTERS_reg_7_30_inst : DLH_X1 port map( G => n11949, D => N3825, Q 
                           => NEXT_REGISTERS_7_30_port);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => N1588, CK => CLK, Q => 
                           n10347, QN => n482_port);
   NEXT_REGISTERS_reg_7_29_inst : DLH_X1 port map( G => n11949, D => N3824, Q 
                           => NEXT_REGISTERS_7_29_port);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => N1587, CK => CLK, Q => 
                           n10345, QN => n483_port);
   NEXT_REGISTERS_reg_7_28_inst : DLH_X1 port map( G => n11949, D => N3823, Q 
                           => NEXT_REGISTERS_7_28_port);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => N1586, CK => CLK, Q => 
                           n10343, QN => n484_port);
   NEXT_REGISTERS_reg_7_27_inst : DLH_X1 port map( G => n11949, D => N3822, Q 
                           => NEXT_REGISTERS_7_27_port);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => N1585, CK => CLK, Q => 
                           n10341, QN => n485_port);
   NEXT_REGISTERS_reg_7_26_inst : DLH_X1 port map( G => n11949, D => N3821, Q 
                           => NEXT_REGISTERS_7_26_port);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => N1584, CK => CLK, Q => 
                           n10339, QN => n486_port);
   NEXT_REGISTERS_reg_7_25_inst : DLH_X1 port map( G => n11949, D => N3820, Q 
                           => NEXT_REGISTERS_7_25_port);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => N1583, CK => CLK, Q => 
                           n10337, QN => n487_port);
   NEXT_REGISTERS_reg_7_24_inst : DLH_X1 port map( G => n11949, D => N3819, Q 
                           => NEXT_REGISTERS_7_24_port);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => N1582, CK => CLK, Q => 
                           n10335, QN => n488_port);
   NEXT_REGISTERS_reg_7_23_inst : DLH_X1 port map( G => n11949, D => N3818, Q 
                           => NEXT_REGISTERS_7_23_port);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => N1581, CK => CLK, Q => 
                           n10333, QN => n489_port);
   NEXT_REGISTERS_reg_7_22_inst : DLH_X1 port map( G => n11949, D => N3817, Q 
                           => NEXT_REGISTERS_7_22_port);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => N1580, CK => CLK, Q => 
                           n10331, QN => n490_port);
   NEXT_REGISTERS_reg_7_21_inst : DLH_X1 port map( G => n11949, D => N3816, Q 
                           => NEXT_REGISTERS_7_21_port);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => N1579, CK => CLK, Q => 
                           n10329, QN => n491_port);
   NEXT_REGISTERS_reg_7_20_inst : DLH_X1 port map( G => n11949, D => N3815, Q 
                           => NEXT_REGISTERS_7_20_port);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => N1578, CK => CLK, Q => 
                           n10327, QN => n492_port);
   NEXT_REGISTERS_reg_7_19_inst : DLH_X1 port map( G => n11950, D => N3814, Q 
                           => NEXT_REGISTERS_7_19_port);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => N1577, CK => CLK, Q => 
                           n10325, QN => n493_port);
   NEXT_REGISTERS_reg_7_18_inst : DLH_X1 port map( G => n11950, D => N3813, Q 
                           => NEXT_REGISTERS_7_18_port);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => N1576, CK => CLK, Q => 
                           n10323, QN => n494_port);
   NEXT_REGISTERS_reg_7_17_inst : DLH_X1 port map( G => n11950, D => N3812, Q 
                           => NEXT_REGISTERS_7_17_port);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => N1575, CK => CLK, Q => 
                           n10321, QN => n495_port);
   NEXT_REGISTERS_reg_7_16_inst : DLH_X1 port map( G => n11950, D => N3811, Q 
                           => NEXT_REGISTERS_7_16_port);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => N1574, CK => CLK, Q => 
                           n10319, QN => n496_port);
   NEXT_REGISTERS_reg_7_15_inst : DLH_X1 port map( G => n11950, D => N3810, Q 
                           => NEXT_REGISTERS_7_15_port);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => N1573, CK => CLK, Q => 
                           n10317, QN => n497_port);
   NEXT_REGISTERS_reg_7_14_inst : DLH_X1 port map( G => n11950, D => N3809, Q 
                           => NEXT_REGISTERS_7_14_port);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => N1572, CK => CLK, Q => 
                           n10315, QN => n498_port);
   NEXT_REGISTERS_reg_7_13_inst : DLH_X1 port map( G => n11950, D => N3808, Q 
                           => NEXT_REGISTERS_7_13_port);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => N1571, CK => CLK, Q => 
                           n10313, QN => n499_port);
   NEXT_REGISTERS_reg_7_12_inst : DLH_X1 port map( G => n11950, D => N3807, Q 
                           => NEXT_REGISTERS_7_12_port);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => N1570, CK => CLK, Q => 
                           n10311, QN => n500_port);
   NEXT_REGISTERS_reg_7_11_inst : DLH_X1 port map( G => n11950, D => N3806, Q 
                           => NEXT_REGISTERS_7_11_port);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => N1569, CK => CLK, Q => 
                           n10309, QN => n501_port);
   NEXT_REGISTERS_reg_7_10_inst : DLH_X1 port map( G => n11950, D => N3805, Q 
                           => NEXT_REGISTERS_7_10_port);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => N1568, CK => CLK, Q => 
                           n10307, QN => n502_port);
   NEXT_REGISTERS_reg_7_9_inst : DLH_X1 port map( G => n11950, D => N3804, Q =>
                           NEXT_REGISTERS_7_9_port);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => N1567, CK => CLK, Q => n10305
                           , QN => n503_port);
   NEXT_REGISTERS_reg_7_8_inst : DLH_X1 port map( G => n11951, D => N3803, Q =>
                           NEXT_REGISTERS_7_8_port);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => N1566, CK => CLK, Q => n10303
                           , QN => n504_port);
   NEXT_REGISTERS_reg_7_7_inst : DLH_X1 port map( G => n11951, D => N3802, Q =>
                           NEXT_REGISTERS_7_7_port);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => N1565, CK => CLK, Q => n10301
                           , QN => n505_port);
   NEXT_REGISTERS_reg_7_6_inst : DLH_X1 port map( G => n11951, D => N3801, Q =>
                           NEXT_REGISTERS_7_6_port);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => N1564, CK => CLK, Q => n10299
                           , QN => n506_port);
   NEXT_REGISTERS_reg_7_5_inst : DLH_X1 port map( G => n11951, D => N3800, Q =>
                           NEXT_REGISTERS_7_5_port);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => N1563, CK => CLK, Q => n10297
                           , QN => n507_port);
   NEXT_REGISTERS_reg_7_4_inst : DLH_X1 port map( G => n11951, D => N3799, Q =>
                           NEXT_REGISTERS_7_4_port);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => N1562, CK => CLK, Q => n10295
                           , QN => n508_port);
   NEXT_REGISTERS_reg_7_3_inst : DLH_X1 port map( G => n11951, D => N3798, Q =>
                           NEXT_REGISTERS_7_3_port);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => N1561, CK => CLK, Q => n10293
                           , QN => n509_port);
   NEXT_REGISTERS_reg_7_2_inst : DLH_X1 port map( G => n11951, D => N3797, Q =>
                           NEXT_REGISTERS_7_2_port);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => N1560, CK => CLK, Q => n10291
                           , QN => n510_port);
   NEXT_REGISTERS_reg_7_1_inst : DLH_X1 port map( G => n11951, D => N3796, Q =>
                           NEXT_REGISTERS_7_1_port);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => N1559, CK => CLK, Q => n10289
                           , QN => n511_port);
   NEXT_REGISTERS_reg_7_0_inst : DLH_X1 port map( G => n11951, D => N3795, Q =>
                           NEXT_REGISTERS_7_0_port);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => N1558, CK => CLK, Q => n10287
                           , QN => n512_port);
   NEXT_REGISTERS_reg_8_63_inst : DLH_X1 port map( G => n11955, D => N3793, Q 
                           => NEXT_REGISTERS_8_63_port);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => N1557, CK => CLK, Q => 
                           n10094, QN => n513_port);
   NEXT_REGISTERS_reg_8_62_inst : DLH_X1 port map( G => n11955, D => N3792, Q 
                           => NEXT_REGISTERS_8_62_port);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => N1556, CK => CLK, Q => 
                           n10092, QN => n514_port);
   NEXT_REGISTERS_reg_8_61_inst : DLH_X1 port map( G => n11955, D => N3791, Q 
                           => NEXT_REGISTERS_8_61_port);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => N1555, CK => CLK, Q => 
                           n10090, QN => n515_port);
   NEXT_REGISTERS_reg_8_60_inst : DLH_X1 port map( G => n11955, D => N3790, Q 
                           => NEXT_REGISTERS_8_60_port);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => N1554, CK => CLK, Q => 
                           n10088, QN => n516_port);
   NEXT_REGISTERS_reg_8_59_inst : DLH_X1 port map( G => n11955, D => N3789, Q 
                           => NEXT_REGISTERS_8_59_port);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => N1553, CK => CLK, Q => 
                           n10086, QN => n517_port);
   NEXT_REGISTERS_reg_8_58_inst : DLH_X1 port map( G => n11955, D => N3788, Q 
                           => NEXT_REGISTERS_8_58_port);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => N1552, CK => CLK, Q => 
                           n10084, QN => n518_port);
   NEXT_REGISTERS_reg_8_57_inst : DLH_X1 port map( G => n11955, D => N3787, Q 
                           => NEXT_REGISTERS_8_57_port);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => N1551, CK => CLK, Q => 
                           n10082, QN => n519_port);
   NEXT_REGISTERS_reg_8_56_inst : DLH_X1 port map( G => n11955, D => N3786, Q 
                           => NEXT_REGISTERS_8_56_port);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => N1550, CK => CLK, Q => 
                           n10080, QN => n520_port);
   NEXT_REGISTERS_reg_8_55_inst : DLH_X1 port map( G => n11955, D => N3785, Q 
                           => NEXT_REGISTERS_8_55_port);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => N1549, CK => CLK, Q => 
                           n10078, QN => n521_port);
   NEXT_REGISTERS_reg_8_54_inst : DLH_X1 port map( G => n11955, D => N3784, Q 
                           => NEXT_REGISTERS_8_54_port);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => N1548, CK => CLK, Q => 
                           n10076, QN => n522_port);
   NEXT_REGISTERS_reg_8_53_inst : DLH_X1 port map( G => n11955, D => N3783, Q 
                           => NEXT_REGISTERS_8_53_port);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => N1547, CK => CLK, Q => 
                           n10074, QN => n523_port);
   NEXT_REGISTERS_reg_8_52_inst : DLH_X1 port map( G => n11956, D => N3782, Q 
                           => NEXT_REGISTERS_8_52_port);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => N1546, CK => CLK, Q => 
                           n10072, QN => n524_port);
   NEXT_REGISTERS_reg_8_51_inst : DLH_X1 port map( G => n11956, D => N3781, Q 
                           => NEXT_REGISTERS_8_51_port);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => N1545, CK => CLK, Q => 
                           n10070, QN => n525_port);
   NEXT_REGISTERS_reg_8_50_inst : DLH_X1 port map( G => n11956, D => N3780, Q 
                           => NEXT_REGISTERS_8_50_port);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => N1544, CK => CLK, Q => 
                           n10068, QN => n526_port);
   NEXT_REGISTERS_reg_8_49_inst : DLH_X1 port map( G => n11956, D => N3779, Q 
                           => NEXT_REGISTERS_8_49_port);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => N1543, CK => CLK, Q => 
                           n10066, QN => n527_port);
   NEXT_REGISTERS_reg_8_48_inst : DLH_X1 port map( G => n11956, D => N3778, Q 
                           => NEXT_REGISTERS_8_48_port);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => N1542, CK => CLK, Q => 
                           n10064, QN => n528_port);
   NEXT_REGISTERS_reg_8_47_inst : DLH_X1 port map( G => n11956, D => N3777, Q 
                           => NEXT_REGISTERS_8_47_port);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => N1541, CK => CLK, Q => 
                           n10062, QN => n529_port);
   NEXT_REGISTERS_reg_8_46_inst : DLH_X1 port map( G => n11956, D => N3776, Q 
                           => NEXT_REGISTERS_8_46_port);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => N1540, CK => CLK, Q => 
                           n10060, QN => n530_port);
   NEXT_REGISTERS_reg_8_45_inst : DLH_X1 port map( G => n11956, D => N3775, Q 
                           => NEXT_REGISTERS_8_45_port);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => N1539, CK => CLK, Q => 
                           n10058, QN => n531_port);
   NEXT_REGISTERS_reg_8_44_inst : DLH_X1 port map( G => n11956, D => N3774, Q 
                           => NEXT_REGISTERS_8_44_port);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => N1538, CK => CLK, Q => 
                           n10056, QN => n532_port);
   NEXT_REGISTERS_reg_8_43_inst : DLH_X1 port map( G => n11956, D => N3773, Q 
                           => NEXT_REGISTERS_8_43_port);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => N1537, CK => CLK, Q => 
                           n10054, QN => n533_port);
   NEXT_REGISTERS_reg_8_42_inst : DLH_X1 port map( G => n11956, D => N3772, Q 
                           => NEXT_REGISTERS_8_42_port);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => N1536, CK => CLK, Q => 
                           n10052, QN => n534_port);
   NEXT_REGISTERS_reg_8_41_inst : DLH_X1 port map( G => n11957, D => N3771, Q 
                           => NEXT_REGISTERS_8_41_port);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => N1535, CK => CLK, Q => 
                           n10050, QN => n535_port);
   NEXT_REGISTERS_reg_8_40_inst : DLH_X1 port map( G => n11957, D => N3770, Q 
                           => NEXT_REGISTERS_8_40_port);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => N1534, CK => CLK, Q => 
                           n10048, QN => n536_port);
   NEXT_REGISTERS_reg_8_39_inst : DLH_X1 port map( G => n11957, D => N3769, Q 
                           => NEXT_REGISTERS_8_39_port);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => N1533, CK => CLK, Q => 
                           n10046, QN => n537_port);
   NEXT_REGISTERS_reg_8_38_inst : DLH_X1 port map( G => n11957, D => N3768, Q 
                           => NEXT_REGISTERS_8_38_port);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => N1532, CK => CLK, Q => 
                           n10044, QN => n538_port);
   NEXT_REGISTERS_reg_8_37_inst : DLH_X1 port map( G => n11957, D => N3767, Q 
                           => NEXT_REGISTERS_8_37_port);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => N1531, CK => CLK, Q => 
                           n10042, QN => n539_port);
   NEXT_REGISTERS_reg_8_36_inst : DLH_X1 port map( G => n11957, D => N3766, Q 
                           => NEXT_REGISTERS_8_36_port);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => N1530, CK => CLK, Q => 
                           n10040, QN => n540_port);
   NEXT_REGISTERS_reg_8_35_inst : DLH_X1 port map( G => n11957, D => N3765, Q 
                           => NEXT_REGISTERS_8_35_port);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => N1529, CK => CLK, Q => 
                           n10038, QN => n541_port);
   NEXT_REGISTERS_reg_8_34_inst : DLH_X1 port map( G => n11957, D => N3764, Q 
                           => NEXT_REGISTERS_8_34_port);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => N1528, CK => CLK, Q => 
                           n10036, QN => n542_port);
   NEXT_REGISTERS_reg_8_33_inst : DLH_X1 port map( G => n11957, D => N3763, Q 
                           => NEXT_REGISTERS_8_33_port);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => N1527, CK => CLK, Q => 
                           n10034, QN => n543_port);
   NEXT_REGISTERS_reg_8_32_inst : DLH_X1 port map( G => n11957, D => N3762, Q 
                           => NEXT_REGISTERS_8_32_port);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => N1526, CK => CLK, Q => 
                           n10032, QN => n544_port);
   NEXT_REGISTERS_reg_8_31_inst : DLH_X1 port map( G => n11957, D => N3761, Q 
                           => NEXT_REGISTERS_8_31_port);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => N1525, CK => CLK, Q => 
                           n10030, QN => n545_port);
   NEXT_REGISTERS_reg_8_30_inst : DLH_X1 port map( G => n11958, D => N3760, Q 
                           => NEXT_REGISTERS_8_30_port);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => N1524, CK => CLK, Q => 
                           n10028, QN => n546_port);
   NEXT_REGISTERS_reg_8_29_inst : DLH_X1 port map( G => n11958, D => N3759, Q 
                           => NEXT_REGISTERS_8_29_port);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => N1523, CK => CLK, Q => 
                           n10026, QN => n547_port);
   NEXT_REGISTERS_reg_8_28_inst : DLH_X1 port map( G => n11958, D => N3758, Q 
                           => NEXT_REGISTERS_8_28_port);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => N1522, CK => CLK, Q => 
                           n10024, QN => n548_port);
   NEXT_REGISTERS_reg_8_27_inst : DLH_X1 port map( G => n11958, D => N3757, Q 
                           => NEXT_REGISTERS_8_27_port);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => N1521, CK => CLK, Q => 
                           n10022, QN => n549_port);
   NEXT_REGISTERS_reg_8_26_inst : DLH_X1 port map( G => n11958, D => N3756, Q 
                           => NEXT_REGISTERS_8_26_port);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => N1520, CK => CLK, Q => 
                           n10020, QN => n550_port);
   NEXT_REGISTERS_reg_8_25_inst : DLH_X1 port map( G => n11958, D => N3755, Q 
                           => NEXT_REGISTERS_8_25_port);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => N1519, CK => CLK, Q => 
                           n10018, QN => n551_port);
   NEXT_REGISTERS_reg_8_24_inst : DLH_X1 port map( G => n11958, D => N3754, Q 
                           => NEXT_REGISTERS_8_24_port);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => N1518, CK => CLK, Q => 
                           n10016, QN => n552_port);
   NEXT_REGISTERS_reg_8_23_inst : DLH_X1 port map( G => n11958, D => N3753, Q 
                           => NEXT_REGISTERS_8_23_port);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => N1517, CK => CLK, Q => 
                           n10014, QN => n553_port);
   NEXT_REGISTERS_reg_8_22_inst : DLH_X1 port map( G => n11958, D => N3752, Q 
                           => NEXT_REGISTERS_8_22_port);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => N1516, CK => CLK, Q => 
                           n10012, QN => n554_port);
   NEXT_REGISTERS_reg_8_21_inst : DLH_X1 port map( G => n11958, D => N3751, Q 
                           => NEXT_REGISTERS_8_21_port);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => N1515, CK => CLK, Q => 
                           n10010, QN => n555_port);
   NEXT_REGISTERS_reg_8_20_inst : DLH_X1 port map( G => n11958, D => N3750, Q 
                           => NEXT_REGISTERS_8_20_port);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => N1514, CK => CLK, Q => 
                           n10008, QN => n556_port);
   NEXT_REGISTERS_reg_8_19_inst : DLH_X1 port map( G => n11959, D => N3749, Q 
                           => NEXT_REGISTERS_8_19_port);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => N1513, CK => CLK, Q => 
                           n10006, QN => n557_port);
   NEXT_REGISTERS_reg_8_18_inst : DLH_X1 port map( G => n11959, D => N3748, Q 
                           => NEXT_REGISTERS_8_18_port);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => N1512, CK => CLK, Q => 
                           n10004, QN => n558_port);
   NEXT_REGISTERS_reg_8_17_inst : DLH_X1 port map( G => n11959, D => N3747, Q 
                           => NEXT_REGISTERS_8_17_port);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => N1511, CK => CLK, Q => 
                           n10002, QN => n559_port);
   NEXT_REGISTERS_reg_8_16_inst : DLH_X1 port map( G => n11959, D => N3746, Q 
                           => NEXT_REGISTERS_8_16_port);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => N1510, CK => CLK, Q => 
                           n10000, QN => n560_port);
   NEXT_REGISTERS_reg_8_15_inst : DLH_X1 port map( G => n11959, D => N3745, Q 
                           => NEXT_REGISTERS_8_15_port);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => N1509, CK => CLK, Q => n9998
                           , QN => n561_port);
   NEXT_REGISTERS_reg_8_14_inst : DLH_X1 port map( G => n11959, D => N3744, Q 
                           => NEXT_REGISTERS_8_14_port);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => N1508, CK => CLK, Q => n9996
                           , QN => n562_port);
   NEXT_REGISTERS_reg_8_13_inst : DLH_X1 port map( G => n11959, D => N3743, Q 
                           => NEXT_REGISTERS_8_13_port);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => N1507, CK => CLK, Q => n9994
                           , QN => n563_port);
   NEXT_REGISTERS_reg_8_12_inst : DLH_X1 port map( G => n11959, D => N3742, Q 
                           => NEXT_REGISTERS_8_12_port);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => N1506, CK => CLK, Q => n9992
                           , QN => n564_port);
   NEXT_REGISTERS_reg_8_11_inst : DLH_X1 port map( G => n11959, D => N3741, Q 
                           => NEXT_REGISTERS_8_11_port);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => N1505, CK => CLK, Q => n9990
                           , QN => n565_port);
   NEXT_REGISTERS_reg_8_10_inst : DLH_X1 port map( G => n11959, D => N3740, Q 
                           => NEXT_REGISTERS_8_10_port);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => N1504, CK => CLK, Q => n9988
                           , QN => n566_port);
   NEXT_REGISTERS_reg_8_9_inst : DLH_X1 port map( G => n11959, D => N3739, Q =>
                           NEXT_REGISTERS_8_9_port);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => N1503, CK => CLK, Q => n9986,
                           QN => n567_port);
   NEXT_REGISTERS_reg_8_8_inst : DLH_X1 port map( G => n11960, D => N3738, Q =>
                           NEXT_REGISTERS_8_8_port);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => N1502, CK => CLK, Q => n9984,
                           QN => n568_port);
   NEXT_REGISTERS_reg_8_7_inst : DLH_X1 port map( G => n11960, D => N3737, Q =>
                           NEXT_REGISTERS_8_7_port);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => N1501, CK => CLK, Q => n9982,
                           QN => n569_port);
   NEXT_REGISTERS_reg_8_6_inst : DLH_X1 port map( G => n11960, D => N3736, Q =>
                           NEXT_REGISTERS_8_6_port);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => N1500, CK => CLK, Q => n9980,
                           QN => n570_port);
   NEXT_REGISTERS_reg_8_5_inst : DLH_X1 port map( G => n11960, D => N3735, Q =>
                           NEXT_REGISTERS_8_5_port);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => N1499, CK => CLK, Q => n9978,
                           QN => n571_port);
   NEXT_REGISTERS_reg_8_4_inst : DLH_X1 port map( G => n11960, D => N3734, Q =>
                           NEXT_REGISTERS_8_4_port);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => N1498, CK => CLK, Q => n9976,
                           QN => n572_port);
   NEXT_REGISTERS_reg_8_3_inst : DLH_X1 port map( G => n11960, D => N3733, Q =>
                           NEXT_REGISTERS_8_3_port);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => N1497, CK => CLK, Q => n9974,
                           QN => n573_port);
   NEXT_REGISTERS_reg_8_2_inst : DLH_X1 port map( G => n11960, D => N3732, Q =>
                           NEXT_REGISTERS_8_2_port);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => N1496, CK => CLK, Q => n9972,
                           QN => n574_port);
   NEXT_REGISTERS_reg_8_1_inst : DLH_X1 port map( G => n11960, D => N3731, Q =>
                           NEXT_REGISTERS_8_1_port);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => N1495, CK => CLK, Q => n9970,
                           QN => n575_port);
   NEXT_REGISTERS_reg_8_0_inst : DLH_X1 port map( G => n11960, D => N3730, Q =>
                           NEXT_REGISTERS_8_0_port);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => N1494, CK => CLK, Q => n9968,
                           QN => n576_port);
   NEXT_REGISTERS_reg_9_63_inst : DLH_X1 port map( G => n11964, D => N3728, Q 
                           => NEXT_REGISTERS_9_63_port);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => N1493, CK => CLK, Q => 
                           n_1256, QN => n577_port);
   NEXT_REGISTERS_reg_9_62_inst : DLH_X1 port map( G => n11964, D => N3727, Q 
                           => NEXT_REGISTERS_9_62_port);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => N1492, CK => CLK, Q => 
                           n_1257, QN => n578_port);
   NEXT_REGISTERS_reg_9_61_inst : DLH_X1 port map( G => n11964, D => N3726, Q 
                           => NEXT_REGISTERS_9_61_port);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => N1491, CK => CLK, Q => 
                           n_1258, QN => n579_port);
   NEXT_REGISTERS_reg_9_60_inst : DLH_X1 port map( G => n11964, D => N3725, Q 
                           => NEXT_REGISTERS_9_60_port);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => N1490, CK => CLK, Q => 
                           n_1259, QN => n580_port);
   NEXT_REGISTERS_reg_9_59_inst : DLH_X1 port map( G => n11964, D => N3724, Q 
                           => NEXT_REGISTERS_9_59_port);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => N1489, CK => CLK, Q => 
                           n_1260, QN => n581_port);
   NEXT_REGISTERS_reg_9_58_inst : DLH_X1 port map( G => n11964, D => N3723, Q 
                           => NEXT_REGISTERS_9_58_port);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => N1488, CK => CLK, Q => 
                           n_1261, QN => n582_port);
   NEXT_REGISTERS_reg_9_57_inst : DLH_X1 port map( G => n11964, D => N3722, Q 
                           => NEXT_REGISTERS_9_57_port);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => N1487, CK => CLK, Q => 
                           n_1262, QN => n583_port);
   NEXT_REGISTERS_reg_9_56_inst : DLH_X1 port map( G => n11964, D => N3721, Q 
                           => NEXT_REGISTERS_9_56_port);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => N1486, CK => CLK, Q => 
                           n_1263, QN => n584_port);
   NEXT_REGISTERS_reg_9_55_inst : DLH_X1 port map( G => n11964, D => N3720, Q 
                           => NEXT_REGISTERS_9_55_port);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => N1485, CK => CLK, Q => 
                           n_1264, QN => n585_port);
   NEXT_REGISTERS_reg_9_54_inst : DLH_X1 port map( G => n11964, D => N3719, Q 
                           => NEXT_REGISTERS_9_54_port);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => N1484, CK => CLK, Q => 
                           n_1265, QN => n586_port);
   NEXT_REGISTERS_reg_9_53_inst : DLH_X1 port map( G => n11964, D => N3718, Q 
                           => NEXT_REGISTERS_9_53_port);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => N1483, CK => CLK, Q => 
                           n_1266, QN => n587_port);
   NEXT_REGISTERS_reg_9_52_inst : DLH_X1 port map( G => n11965, D => N3717, Q 
                           => NEXT_REGISTERS_9_52_port);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => N1482, CK => CLK, Q => 
                           n_1267, QN => n588_port);
   NEXT_REGISTERS_reg_9_51_inst : DLH_X1 port map( G => n11965, D => N3716, Q 
                           => NEXT_REGISTERS_9_51_port);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => N1481, CK => CLK, Q => 
                           n_1268, QN => n589_port);
   NEXT_REGISTERS_reg_9_50_inst : DLH_X1 port map( G => n11965, D => N3715, Q 
                           => NEXT_REGISTERS_9_50_port);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => N1480, CK => CLK, Q => 
                           n_1269, QN => n590_port);
   NEXT_REGISTERS_reg_9_49_inst : DLH_X1 port map( G => n11965, D => N3714, Q 
                           => NEXT_REGISTERS_9_49_port);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => N1479, CK => CLK, Q => 
                           n_1270, QN => n591_port);
   NEXT_REGISTERS_reg_9_48_inst : DLH_X1 port map( G => n11965, D => N3713, Q 
                           => NEXT_REGISTERS_9_48_port);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => N1478, CK => CLK, Q => 
                           n_1271, QN => n592_port);
   NEXT_REGISTERS_reg_9_47_inst : DLH_X1 port map( G => n11965, D => N3712, Q 
                           => NEXT_REGISTERS_9_47_port);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => N1477, CK => CLK, Q => 
                           n_1272, QN => n593_port);
   NEXT_REGISTERS_reg_9_46_inst : DLH_X1 port map( G => n11965, D => N3711, Q 
                           => NEXT_REGISTERS_9_46_port);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => N1476, CK => CLK, Q => 
                           n_1273, QN => n594_port);
   NEXT_REGISTERS_reg_9_45_inst : DLH_X1 port map( G => n11965, D => N3710, Q 
                           => NEXT_REGISTERS_9_45_port);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => N1475, CK => CLK, Q => 
                           n_1274, QN => n595_port);
   NEXT_REGISTERS_reg_9_44_inst : DLH_X1 port map( G => n11965, D => N3709, Q 
                           => NEXT_REGISTERS_9_44_port);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => N1474, CK => CLK, Q => 
                           n_1275, QN => n596_port);
   NEXT_REGISTERS_reg_9_43_inst : DLH_X1 port map( G => n11965, D => N3708, Q 
                           => NEXT_REGISTERS_9_43_port);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => N1473, CK => CLK, Q => 
                           n_1276, QN => n597_port);
   NEXT_REGISTERS_reg_9_42_inst : DLH_X1 port map( G => n11965, D => N3707, Q 
                           => NEXT_REGISTERS_9_42_port);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => N1472, CK => CLK, Q => 
                           n_1277, QN => n598_port);
   NEXT_REGISTERS_reg_9_41_inst : DLH_X1 port map( G => n11966, D => N3706, Q 
                           => NEXT_REGISTERS_9_41_port);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => N1471, CK => CLK, Q => 
                           n_1278, QN => n599_port);
   NEXT_REGISTERS_reg_9_40_inst : DLH_X1 port map( G => n11966, D => N3705, Q 
                           => NEXT_REGISTERS_9_40_port);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => N1470, CK => CLK, Q => 
                           n_1279, QN => n600_port);
   NEXT_REGISTERS_reg_9_39_inst : DLH_X1 port map( G => n11966, D => N3704, Q 
                           => NEXT_REGISTERS_9_39_port);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => N1469, CK => CLK, Q => 
                           n_1280, QN => n601_port);
   NEXT_REGISTERS_reg_9_38_inst : DLH_X1 port map( G => n11966, D => N3703, Q 
                           => NEXT_REGISTERS_9_38_port);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => N1468, CK => CLK, Q => 
                           n_1281, QN => n602_port);
   NEXT_REGISTERS_reg_9_37_inst : DLH_X1 port map( G => n11966, D => N3702, Q 
                           => NEXT_REGISTERS_9_37_port);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => N1467, CK => CLK, Q => 
                           n_1282, QN => n603_port);
   NEXT_REGISTERS_reg_9_36_inst : DLH_X1 port map( G => n11966, D => N3701, Q 
                           => NEXT_REGISTERS_9_36_port);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => N1466, CK => CLK, Q => 
                           n_1283, QN => n604_port);
   NEXT_REGISTERS_reg_9_35_inst : DLH_X1 port map( G => n11966, D => N3700, Q 
                           => NEXT_REGISTERS_9_35_port);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => N1465, CK => CLK, Q => 
                           n_1284, QN => n605_port);
   NEXT_REGISTERS_reg_9_34_inst : DLH_X1 port map( G => n11966, D => N3699, Q 
                           => NEXT_REGISTERS_9_34_port);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => N1464, CK => CLK, Q => 
                           n_1285, QN => n606_port);
   NEXT_REGISTERS_reg_9_33_inst : DLH_X1 port map( G => n11966, D => N3698, Q 
                           => NEXT_REGISTERS_9_33_port);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => N1463, CK => CLK, Q => 
                           n_1286, QN => n607_port);
   NEXT_REGISTERS_reg_9_32_inst : DLH_X1 port map( G => n11966, D => N3697, Q 
                           => NEXT_REGISTERS_9_32_port);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => N1462, CK => CLK, Q => 
                           n_1287, QN => n608_port);
   NEXT_REGISTERS_reg_9_31_inst : DLH_X1 port map( G => n11966, D => N3696, Q 
                           => NEXT_REGISTERS_9_31_port);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => N1461, CK => CLK, Q => 
                           n_1288, QN => n609_port);
   NEXT_REGISTERS_reg_9_30_inst : DLH_X1 port map( G => n11967, D => N3695, Q 
                           => NEXT_REGISTERS_9_30_port);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => N1460, CK => CLK, Q => 
                           n_1289, QN => n610_port);
   NEXT_REGISTERS_reg_9_29_inst : DLH_X1 port map( G => n11967, D => N3694, Q 
                           => NEXT_REGISTERS_9_29_port);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => N1459, CK => CLK, Q => 
                           n_1290, QN => n611_port);
   NEXT_REGISTERS_reg_9_28_inst : DLH_X1 port map( G => n11967, D => N3693, Q 
                           => NEXT_REGISTERS_9_28_port);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => N1458, CK => CLK, Q => 
                           n_1291, QN => n612_port);
   NEXT_REGISTERS_reg_9_27_inst : DLH_X1 port map( G => n11967, D => N3692, Q 
                           => NEXT_REGISTERS_9_27_port);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => N1457, CK => CLK, Q => 
                           n_1292, QN => n613_port);
   NEXT_REGISTERS_reg_9_26_inst : DLH_X1 port map( G => n11967, D => N3691, Q 
                           => NEXT_REGISTERS_9_26_port);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => N1456, CK => CLK, Q => 
                           n_1293, QN => n614_port);
   NEXT_REGISTERS_reg_9_25_inst : DLH_X1 port map( G => n11967, D => N3690, Q 
                           => NEXT_REGISTERS_9_25_port);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => N1455, CK => CLK, Q => 
                           n_1294, QN => n615_port);
   NEXT_REGISTERS_reg_9_24_inst : DLH_X1 port map( G => n11967, D => N3689, Q 
                           => NEXT_REGISTERS_9_24_port);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => N1454, CK => CLK, Q => 
                           n_1295, QN => n616_port);
   NEXT_REGISTERS_reg_9_23_inst : DLH_X1 port map( G => n11967, D => N3688, Q 
                           => NEXT_REGISTERS_9_23_port);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => N1453, CK => CLK, Q => 
                           n_1296, QN => n617_port);
   NEXT_REGISTERS_reg_9_22_inst : DLH_X1 port map( G => n11967, D => N3687, Q 
                           => NEXT_REGISTERS_9_22_port);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => N1452, CK => CLK, Q => 
                           n_1297, QN => n618_port);
   NEXT_REGISTERS_reg_9_21_inst : DLH_X1 port map( G => n11967, D => N3686, Q 
                           => NEXT_REGISTERS_9_21_port);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => N1451, CK => CLK, Q => 
                           n_1298, QN => n619_port);
   NEXT_REGISTERS_reg_9_20_inst : DLH_X1 port map( G => n11967, D => N3685, Q 
                           => NEXT_REGISTERS_9_20_port);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => N1450, CK => CLK, Q => 
                           n_1299, QN => n620_port);
   NEXT_REGISTERS_reg_9_19_inst : DLH_X1 port map( G => n11968, D => N3684, Q 
                           => NEXT_REGISTERS_9_19_port);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => N1449, CK => CLK, Q => 
                           n_1300, QN => n621_port);
   NEXT_REGISTERS_reg_9_18_inst : DLH_X1 port map( G => n11968, D => N3683, Q 
                           => NEXT_REGISTERS_9_18_port);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => N1448, CK => CLK, Q => 
                           n_1301, QN => n622_port);
   NEXT_REGISTERS_reg_9_17_inst : DLH_X1 port map( G => n11968, D => N3682, Q 
                           => NEXT_REGISTERS_9_17_port);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => N1447, CK => CLK, Q => 
                           n_1302, QN => n623_port);
   NEXT_REGISTERS_reg_9_16_inst : DLH_X1 port map( G => n11968, D => N3681, Q 
                           => NEXT_REGISTERS_9_16_port);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => N1446, CK => CLK, Q => 
                           n_1303, QN => n624_port);
   NEXT_REGISTERS_reg_9_15_inst : DLH_X1 port map( G => n11968, D => N3680, Q 
                           => NEXT_REGISTERS_9_15_port);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => N1445, CK => CLK, Q => 
                           n_1304, QN => n625_port);
   NEXT_REGISTERS_reg_9_14_inst : DLH_X1 port map( G => n11968, D => N3679, Q 
                           => NEXT_REGISTERS_9_14_port);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => N1444, CK => CLK, Q => 
                           n_1305, QN => n626_port);
   NEXT_REGISTERS_reg_9_13_inst : DLH_X1 port map( G => n11968, D => N3678, Q 
                           => NEXT_REGISTERS_9_13_port);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => N1443, CK => CLK, Q => 
                           n_1306, QN => n627_port);
   NEXT_REGISTERS_reg_9_12_inst : DLH_X1 port map( G => n11968, D => N3677, Q 
                           => NEXT_REGISTERS_9_12_port);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => N1442, CK => CLK, Q => 
                           n_1307, QN => n628_port);
   NEXT_REGISTERS_reg_9_11_inst : DLH_X1 port map( G => n11968, D => N3676, Q 
                           => NEXT_REGISTERS_9_11_port);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => N1441, CK => CLK, Q => 
                           n_1308, QN => n629_port);
   NEXT_REGISTERS_reg_9_10_inst : DLH_X1 port map( G => n11968, D => N3675, Q 
                           => NEXT_REGISTERS_9_10_port);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => N1440, CK => CLK, Q => 
                           n_1309, QN => n630_port);
   NEXT_REGISTERS_reg_9_9_inst : DLH_X1 port map( G => n11968, D => N3674, Q =>
                           NEXT_REGISTERS_9_9_port);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => N1439, CK => CLK, Q => n_1310
                           , QN => n631_port);
   NEXT_REGISTERS_reg_9_8_inst : DLH_X1 port map( G => n11969, D => N3673, Q =>
                           NEXT_REGISTERS_9_8_port);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => N1438, CK => CLK, Q => n_1311
                           , QN => n632_port);
   NEXT_REGISTERS_reg_9_7_inst : DLH_X1 port map( G => n11969, D => N3672, Q =>
                           NEXT_REGISTERS_9_7_port);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => N1437, CK => CLK, Q => n_1312
                           , QN => n633_port);
   NEXT_REGISTERS_reg_9_6_inst : DLH_X1 port map( G => n11969, D => N3671, Q =>
                           NEXT_REGISTERS_9_6_port);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => N1436, CK => CLK, Q => n_1313
                           , QN => n634_port);
   NEXT_REGISTERS_reg_9_5_inst : DLH_X1 port map( G => n11969, D => N3670, Q =>
                           NEXT_REGISTERS_9_5_port);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => N1435, CK => CLK, Q => n_1314
                           , QN => n635_port);
   NEXT_REGISTERS_reg_9_4_inst : DLH_X1 port map( G => n11969, D => N3669, Q =>
                           NEXT_REGISTERS_9_4_port);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => N1434, CK => CLK, Q => n_1315
                           , QN => n636_port);
   NEXT_REGISTERS_reg_9_3_inst : DLH_X1 port map( G => n11969, D => N3668, Q =>
                           NEXT_REGISTERS_9_3_port);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => N1433, CK => CLK, Q => n_1316
                           , QN => n637_port);
   NEXT_REGISTERS_reg_9_2_inst : DLH_X1 port map( G => n11969, D => N3667, Q =>
                           NEXT_REGISTERS_9_2_port);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => N1432, CK => CLK, Q => n_1317
                           , QN => n638_port);
   NEXT_REGISTERS_reg_9_1_inst : DLH_X1 port map( G => n11969, D => N3666, Q =>
                           NEXT_REGISTERS_9_1_port);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => N1431, CK => CLK, Q => n_1318
                           , QN => n639_port);
   NEXT_REGISTERS_reg_9_0_inst : DLH_X1 port map( G => n11969, D => N3665, Q =>
                           NEXT_REGISTERS_9_0_port);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => N1430, CK => CLK, Q => n_1319
                           , QN => n640_port);
   NEXT_REGISTERS_reg_10_63_inst : DLH_X1 port map( G => n11973, D => N3663, Q 
                           => NEXT_REGISTERS_10_63_port);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => N1429, CK => CLK, Q => 
                           n10542, QN => n641_port);
   NEXT_REGISTERS_reg_10_62_inst : DLH_X1 port map( G => n11973, D => N3662, Q 
                           => NEXT_REGISTERS_10_62_port);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => N1428, CK => CLK, Q => 
                           n10540, QN => n642_port);
   NEXT_REGISTERS_reg_10_61_inst : DLH_X1 port map( G => n11973, D => N3661, Q 
                           => NEXT_REGISTERS_10_61_port);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => N1427, CK => CLK, Q => 
                           n10538, QN => n643_port);
   NEXT_REGISTERS_reg_10_60_inst : DLH_X1 port map( G => n11973, D => N3660, Q 
                           => NEXT_REGISTERS_10_60_port);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => N1426, CK => CLK, Q => 
                           n10536, QN => n644_port);
   NEXT_REGISTERS_reg_10_59_inst : DLH_X1 port map( G => n11973, D => N3659, Q 
                           => NEXT_REGISTERS_10_59_port);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => N1425, CK => CLK, Q => 
                           n10534, QN => n645_port);
   NEXT_REGISTERS_reg_10_58_inst : DLH_X1 port map( G => n11973, D => N3658, Q 
                           => NEXT_REGISTERS_10_58_port);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => N1424, CK => CLK, Q => 
                           n10532, QN => n646_port);
   NEXT_REGISTERS_reg_10_57_inst : DLH_X1 port map( G => n11973, D => N3657, Q 
                           => NEXT_REGISTERS_10_57_port);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => N1423, CK => CLK, Q => 
                           n10530, QN => n647_port);
   NEXT_REGISTERS_reg_10_56_inst : DLH_X1 port map( G => n11973, D => N3656, Q 
                           => NEXT_REGISTERS_10_56_port);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => N1422, CK => CLK, Q => 
                           n10528, QN => n648_port);
   NEXT_REGISTERS_reg_10_55_inst : DLH_X1 port map( G => n11973, D => N3655, Q 
                           => NEXT_REGISTERS_10_55_port);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => N1421, CK => CLK, Q => 
                           n10526, QN => n649_port);
   NEXT_REGISTERS_reg_10_54_inst : DLH_X1 port map( G => n11973, D => N3654, Q 
                           => NEXT_REGISTERS_10_54_port);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => N1420, CK => CLK, Q => 
                           n10524, QN => n650_port);
   NEXT_REGISTERS_reg_10_53_inst : DLH_X1 port map( G => n11973, D => N3653, Q 
                           => NEXT_REGISTERS_10_53_port);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => N1419, CK => CLK, Q => 
                           n10522, QN => n651_port);
   NEXT_REGISTERS_reg_10_52_inst : DLH_X1 port map( G => n11974, D => N3652, Q 
                           => NEXT_REGISTERS_10_52_port);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => N1418, CK => CLK, Q => 
                           n10520, QN => n652_port);
   NEXT_REGISTERS_reg_10_51_inst : DLH_X1 port map( G => n11974, D => N3651, Q 
                           => NEXT_REGISTERS_10_51_port);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => N1417, CK => CLK, Q => 
                           n10518, QN => n653_port);
   NEXT_REGISTERS_reg_10_50_inst : DLH_X1 port map( G => n11974, D => N3650, Q 
                           => NEXT_REGISTERS_10_50_port);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => N1416, CK => CLK, Q => 
                           n10516, QN => n654_port);
   NEXT_REGISTERS_reg_10_49_inst : DLH_X1 port map( G => n11974, D => N3649, Q 
                           => NEXT_REGISTERS_10_49_port);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => N1415, CK => CLK, Q => 
                           n10514, QN => n655_port);
   NEXT_REGISTERS_reg_10_48_inst : DLH_X1 port map( G => n11974, D => N3648, Q 
                           => NEXT_REGISTERS_10_48_port);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => N1414, CK => CLK, Q => 
                           n10512, QN => n656_port);
   NEXT_REGISTERS_reg_10_47_inst : DLH_X1 port map( G => n11974, D => N3647, Q 
                           => NEXT_REGISTERS_10_47_port);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => N1413, CK => CLK, Q => 
                           n10510, QN => n657_port);
   NEXT_REGISTERS_reg_10_46_inst : DLH_X1 port map( G => n11974, D => N3646, Q 
                           => NEXT_REGISTERS_10_46_port);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => N1412, CK => CLK, Q => 
                           n10508, QN => n658_port);
   NEXT_REGISTERS_reg_10_45_inst : DLH_X1 port map( G => n11974, D => N3645, Q 
                           => NEXT_REGISTERS_10_45_port);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => N1411, CK => CLK, Q => 
                           n10506, QN => n659_port);
   NEXT_REGISTERS_reg_10_44_inst : DLH_X1 port map( G => n11974, D => N3644, Q 
                           => NEXT_REGISTERS_10_44_port);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => N1410, CK => CLK, Q => 
                           n10504, QN => n660_port);
   NEXT_REGISTERS_reg_10_43_inst : DLH_X1 port map( G => n11974, D => N3643, Q 
                           => NEXT_REGISTERS_10_43_port);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => N1409, CK => CLK, Q => 
                           n10502, QN => n661_port);
   NEXT_REGISTERS_reg_10_42_inst : DLH_X1 port map( G => n11974, D => N3642, Q 
                           => NEXT_REGISTERS_10_42_port);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => N1408, CK => CLK, Q => 
                           n10500, QN => n662_port);
   NEXT_REGISTERS_reg_10_41_inst : DLH_X1 port map( G => n11975, D => N3641, Q 
                           => NEXT_REGISTERS_10_41_port);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => N1407, CK => CLK, Q => 
                           n10498, QN => n663_port);
   NEXT_REGISTERS_reg_10_40_inst : DLH_X1 port map( G => n11975, D => N3640, Q 
                           => NEXT_REGISTERS_10_40_port);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => N1406, CK => CLK, Q => 
                           n10496, QN => n664_port);
   NEXT_REGISTERS_reg_10_39_inst : DLH_X1 port map( G => n11975, D => N3639, Q 
                           => NEXT_REGISTERS_10_39_port);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => N1405, CK => CLK, Q => 
                           n10494, QN => n665_port);
   NEXT_REGISTERS_reg_10_38_inst : DLH_X1 port map( G => n11975, D => N3638, Q 
                           => NEXT_REGISTERS_10_38_port);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => N1404, CK => CLK, Q => 
                           n10492, QN => n666_port);
   NEXT_REGISTERS_reg_10_37_inst : DLH_X1 port map( G => n11975, D => N3637, Q 
                           => NEXT_REGISTERS_10_37_port);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => N1403, CK => CLK, Q => 
                           n10490, QN => n667_port);
   NEXT_REGISTERS_reg_10_36_inst : DLH_X1 port map( G => n11975, D => N3636, Q 
                           => NEXT_REGISTERS_10_36_port);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => N1402, CK => CLK, Q => 
                           n10488, QN => n668_port);
   NEXT_REGISTERS_reg_10_35_inst : DLH_X1 port map( G => n11975, D => N3635, Q 
                           => NEXT_REGISTERS_10_35_port);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => N1401, CK => CLK, Q => 
                           n10486, QN => n669_port);
   NEXT_REGISTERS_reg_10_34_inst : DLH_X1 port map( G => n11975, D => N3634, Q 
                           => NEXT_REGISTERS_10_34_port);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => N1400, CK => CLK, Q => 
                           n10484, QN => n670_port);
   NEXT_REGISTERS_reg_10_33_inst : DLH_X1 port map( G => n11975, D => N3633, Q 
                           => NEXT_REGISTERS_10_33_port);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => N1399, CK => CLK, Q => 
                           n10482, QN => n671_port);
   NEXT_REGISTERS_reg_10_32_inst : DLH_X1 port map( G => n11975, D => N3632, Q 
                           => NEXT_REGISTERS_10_32_port);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => N1398, CK => CLK, Q => 
                           n10480, QN => n672_port);
   NEXT_REGISTERS_reg_10_31_inst : DLH_X1 port map( G => n11975, D => N3631, Q 
                           => NEXT_REGISTERS_10_31_port);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => N1397, CK => CLK, Q => 
                           n10478, QN => n673_port);
   NEXT_REGISTERS_reg_10_30_inst : DLH_X1 port map( G => n11976, D => N3630, Q 
                           => NEXT_REGISTERS_10_30_port);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => N1396, CK => CLK, Q => 
                           n10476, QN => n674_port);
   NEXT_REGISTERS_reg_10_29_inst : DLH_X1 port map( G => n11976, D => N3629, Q 
                           => NEXT_REGISTERS_10_29_port);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => N1395, CK => CLK, Q => 
                           n10474, QN => n675_port);
   NEXT_REGISTERS_reg_10_28_inst : DLH_X1 port map( G => n11976, D => N3628, Q 
                           => NEXT_REGISTERS_10_28_port);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => N1394, CK => CLK, Q => 
                           n10472, QN => n676_port);
   NEXT_REGISTERS_reg_10_27_inst : DLH_X1 port map( G => n11976, D => N3627, Q 
                           => NEXT_REGISTERS_10_27_port);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => N1393, CK => CLK, Q => 
                           n10470, QN => n677_port);
   NEXT_REGISTERS_reg_10_26_inst : DLH_X1 port map( G => n11976, D => N3626, Q 
                           => NEXT_REGISTERS_10_26_port);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => N1392, CK => CLK, Q => 
                           n10468, QN => n678_port);
   NEXT_REGISTERS_reg_10_25_inst : DLH_X1 port map( G => n11976, D => N3625, Q 
                           => NEXT_REGISTERS_10_25_port);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => N1391, CK => CLK, Q => 
                           n10466, QN => n679_port);
   NEXT_REGISTERS_reg_10_24_inst : DLH_X1 port map( G => n11976, D => N3624, Q 
                           => NEXT_REGISTERS_10_24_port);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => N1390, CK => CLK, Q => 
                           n10464, QN => n680_port);
   NEXT_REGISTERS_reg_10_23_inst : DLH_X1 port map( G => n11976, D => N3623, Q 
                           => NEXT_REGISTERS_10_23_port);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => N1389, CK => CLK, Q => 
                           n10462, QN => n681_port);
   NEXT_REGISTERS_reg_10_22_inst : DLH_X1 port map( G => n11976, D => N3622, Q 
                           => NEXT_REGISTERS_10_22_port);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => N1388, CK => CLK, Q => 
                           n10460, QN => n682_port);
   NEXT_REGISTERS_reg_10_21_inst : DLH_X1 port map( G => n11976, D => N3621, Q 
                           => NEXT_REGISTERS_10_21_port);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => N1387, CK => CLK, Q => 
                           n10458, QN => n683_port);
   NEXT_REGISTERS_reg_10_20_inst : DLH_X1 port map( G => n11976, D => N3620, Q 
                           => NEXT_REGISTERS_10_20_port);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => N1386, CK => CLK, Q => 
                           n10456, QN => n684_port);
   NEXT_REGISTERS_reg_10_19_inst : DLH_X1 port map( G => n11977, D => N3619, Q 
                           => NEXT_REGISTERS_10_19_port);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => N1385, CK => CLK, Q => 
                           n10454, QN => n685_port);
   NEXT_REGISTERS_reg_10_18_inst : DLH_X1 port map( G => n11977, D => N3618, Q 
                           => NEXT_REGISTERS_10_18_port);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => N1384, CK => CLK, Q => 
                           n10452, QN => n686_port);
   NEXT_REGISTERS_reg_10_17_inst : DLH_X1 port map( G => n11977, D => N3617, Q 
                           => NEXT_REGISTERS_10_17_port);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => N1383, CK => CLK, Q => 
                           n10450, QN => n687_port);
   NEXT_REGISTERS_reg_10_16_inst : DLH_X1 port map( G => n11977, D => N3616, Q 
                           => NEXT_REGISTERS_10_16_port);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => N1382, CK => CLK, Q => 
                           n10448, QN => n688_port);
   NEXT_REGISTERS_reg_10_15_inst : DLH_X1 port map( G => n11977, D => N3615, Q 
                           => NEXT_REGISTERS_10_15_port);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => N1381, CK => CLK, Q => 
                           n10446, QN => n689_port);
   NEXT_REGISTERS_reg_10_14_inst : DLH_X1 port map( G => n11977, D => N3614, Q 
                           => NEXT_REGISTERS_10_14_port);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => N1380, CK => CLK, Q => 
                           n10444, QN => n690_port);
   NEXT_REGISTERS_reg_10_13_inst : DLH_X1 port map( G => n11977, D => N3613, Q 
                           => NEXT_REGISTERS_10_13_port);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => N1379, CK => CLK, Q => 
                           n10442, QN => n691_port);
   NEXT_REGISTERS_reg_10_12_inst : DLH_X1 port map( G => n11977, D => N3612, Q 
                           => NEXT_REGISTERS_10_12_port);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => N1378, CK => CLK, Q => 
                           n10440, QN => n692_port);
   NEXT_REGISTERS_reg_10_11_inst : DLH_X1 port map( G => n11977, D => N3611, Q 
                           => NEXT_REGISTERS_10_11_port);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => N1377, CK => CLK, Q => 
                           n10438, QN => n693_port);
   NEXT_REGISTERS_reg_10_10_inst : DLH_X1 port map( G => n11977, D => N3610, Q 
                           => NEXT_REGISTERS_10_10_port);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => N1376, CK => CLK, Q => 
                           n10436, QN => n694_port);
   NEXT_REGISTERS_reg_10_9_inst : DLH_X1 port map( G => n11977, D => N3609, Q 
                           => NEXT_REGISTERS_10_9_port);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => N1375, CK => CLK, Q => 
                           n10434, QN => n695_port);
   NEXT_REGISTERS_reg_10_8_inst : DLH_X1 port map( G => n11978, D => N3608, Q 
                           => NEXT_REGISTERS_10_8_port);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => N1374, CK => CLK, Q => 
                           n10432, QN => n696_port);
   NEXT_REGISTERS_reg_10_7_inst : DLH_X1 port map( G => n11978, D => N3607, Q 
                           => NEXT_REGISTERS_10_7_port);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => N1373, CK => CLK, Q => 
                           n10430, QN => n697_port);
   NEXT_REGISTERS_reg_10_6_inst : DLH_X1 port map( G => n11978, D => N3606, Q 
                           => NEXT_REGISTERS_10_6_port);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => N1372, CK => CLK, Q => 
                           n10428, QN => n698_port);
   NEXT_REGISTERS_reg_10_5_inst : DLH_X1 port map( G => n11978, D => N3605, Q 
                           => NEXT_REGISTERS_10_5_port);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => N1371, CK => CLK, Q => 
                           n10426, QN => n699_port);
   NEXT_REGISTERS_reg_10_4_inst : DLH_X1 port map( G => n11978, D => N3604, Q 
                           => NEXT_REGISTERS_10_4_port);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => N1370, CK => CLK, Q => 
                           n10424, QN => n700_port);
   NEXT_REGISTERS_reg_10_3_inst : DLH_X1 port map( G => n11978, D => N3603, Q 
                           => NEXT_REGISTERS_10_3_port);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => N1369, CK => CLK, Q => 
                           n10422, QN => n701_port);
   NEXT_REGISTERS_reg_10_2_inst : DLH_X1 port map( G => n11978, D => N3602, Q 
                           => NEXT_REGISTERS_10_2_port);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => N1368, CK => CLK, Q => 
                           n10420, QN => n702_port);
   NEXT_REGISTERS_reg_10_1_inst : DLH_X1 port map( G => n11978, D => N3601, Q 
                           => NEXT_REGISTERS_10_1_port);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => N1367, CK => CLK, Q => 
                           n10418, QN => n703_port);
   NEXT_REGISTERS_reg_10_0_inst : DLH_X1 port map( G => n11978, D => N3600, Q 
                           => NEXT_REGISTERS_10_0_port);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => N1366, CK => CLK, Q => 
                           n10416, QN => n704_port);
   NEXT_REGISTERS_reg_11_63_inst : DLH_X1 port map( G => n11982, D => N3598, Q 
                           => NEXT_REGISTERS_11_63_port);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => N1365, CK => CLK, Q => 
                           n_1320, QN => n705_port);
   NEXT_REGISTERS_reg_11_62_inst : DLH_X1 port map( G => n11982, D => N3597, Q 
                           => NEXT_REGISTERS_11_62_port);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => N1364, CK => CLK, Q => 
                           n_1321, QN => n706_port);
   NEXT_REGISTERS_reg_11_61_inst : DLH_X1 port map( G => n11982, D => N3596, Q 
                           => NEXT_REGISTERS_11_61_port);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => N1363, CK => CLK, Q => 
                           n_1322, QN => n707_port);
   NEXT_REGISTERS_reg_11_60_inst : DLH_X1 port map( G => n11982, D => N3595, Q 
                           => NEXT_REGISTERS_11_60_port);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => N1362, CK => CLK, Q => 
                           n_1323, QN => n708_port);
   NEXT_REGISTERS_reg_11_59_inst : DLH_X1 port map( G => n11982, D => N3594, Q 
                           => NEXT_REGISTERS_11_59_port);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => N1361, CK => CLK, Q => 
                           n_1324, QN => n709_port);
   NEXT_REGISTERS_reg_11_58_inst : DLH_X1 port map( G => n11982, D => N3593, Q 
                           => NEXT_REGISTERS_11_58_port);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => N1360, CK => CLK, Q => 
                           n_1325, QN => n710_port);
   NEXT_REGISTERS_reg_11_57_inst : DLH_X1 port map( G => n11982, D => N3592, Q 
                           => NEXT_REGISTERS_11_57_port);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => N1359, CK => CLK, Q => 
                           n_1326, QN => n711_port);
   NEXT_REGISTERS_reg_11_56_inst : DLH_X1 port map( G => n11982, D => N3591, Q 
                           => NEXT_REGISTERS_11_56_port);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => N1358, CK => CLK, Q => 
                           n_1327, QN => n712_port);
   NEXT_REGISTERS_reg_11_55_inst : DLH_X1 port map( G => n11982, D => N3590, Q 
                           => NEXT_REGISTERS_11_55_port);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => N1357, CK => CLK, Q => 
                           n_1328, QN => n713_port);
   NEXT_REGISTERS_reg_11_54_inst : DLH_X1 port map( G => n11982, D => N3589, Q 
                           => NEXT_REGISTERS_11_54_port);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => N1356, CK => CLK, Q => 
                           n_1329, QN => n714_port);
   NEXT_REGISTERS_reg_11_53_inst : DLH_X1 port map( G => n11982, D => N3588, Q 
                           => NEXT_REGISTERS_11_53_port);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => N1355, CK => CLK, Q => 
                           n_1330, QN => n715_port);
   NEXT_REGISTERS_reg_11_52_inst : DLH_X1 port map( G => n11983, D => N3587, Q 
                           => NEXT_REGISTERS_11_52_port);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => N1354, CK => CLK, Q => 
                           n_1331, QN => n716_port);
   NEXT_REGISTERS_reg_11_51_inst : DLH_X1 port map( G => n11983, D => N3586, Q 
                           => NEXT_REGISTERS_11_51_port);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => N1353, CK => CLK, Q => 
                           n_1332, QN => n717_port);
   NEXT_REGISTERS_reg_11_50_inst : DLH_X1 port map( G => n11983, D => N3585, Q 
                           => NEXT_REGISTERS_11_50_port);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => N1352, CK => CLK, Q => 
                           n_1333, QN => n718_port);
   NEXT_REGISTERS_reg_11_49_inst : DLH_X1 port map( G => n11983, D => N3584, Q 
                           => NEXT_REGISTERS_11_49_port);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => N1351, CK => CLK, Q => 
                           n_1334, QN => n719_port);
   NEXT_REGISTERS_reg_11_48_inst : DLH_X1 port map( G => n11983, D => N3583, Q 
                           => NEXT_REGISTERS_11_48_port);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => N1350, CK => CLK, Q => 
                           n_1335, QN => n720_port);
   NEXT_REGISTERS_reg_11_47_inst : DLH_X1 port map( G => n11983, D => N3582, Q 
                           => NEXT_REGISTERS_11_47_port);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => N1349, CK => CLK, Q => 
                           n_1336, QN => n721_port);
   NEXT_REGISTERS_reg_11_46_inst : DLH_X1 port map( G => n11983, D => N3581, Q 
                           => NEXT_REGISTERS_11_46_port);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => N1348, CK => CLK, Q => 
                           n_1337, QN => n722_port);
   NEXT_REGISTERS_reg_11_45_inst : DLH_X1 port map( G => n11983, D => N3580, Q 
                           => NEXT_REGISTERS_11_45_port);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => N1347, CK => CLK, Q => 
                           n_1338, QN => n723_port);
   NEXT_REGISTERS_reg_11_44_inst : DLH_X1 port map( G => n11983, D => N3579, Q 
                           => NEXT_REGISTERS_11_44_port);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => N1346, CK => CLK, Q => 
                           n_1339, QN => n724_port);
   NEXT_REGISTERS_reg_11_43_inst : DLH_X1 port map( G => n11983, D => N3578, Q 
                           => NEXT_REGISTERS_11_43_port);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => N1345, CK => CLK, Q => 
                           n_1340, QN => n725_port);
   NEXT_REGISTERS_reg_11_42_inst : DLH_X1 port map( G => n11983, D => N3577, Q 
                           => NEXT_REGISTERS_11_42_port);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => N1344, CK => CLK, Q => 
                           n_1341, QN => n726_port);
   NEXT_REGISTERS_reg_11_41_inst : DLH_X1 port map( G => n11984, D => N3576, Q 
                           => NEXT_REGISTERS_11_41_port);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => N1343, CK => CLK, Q => 
                           n_1342, QN => n727_port);
   NEXT_REGISTERS_reg_11_40_inst : DLH_X1 port map( G => n11984, D => N3575, Q 
                           => NEXT_REGISTERS_11_40_port);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => N1342, CK => CLK, Q => 
                           n_1343, QN => n728_port);
   NEXT_REGISTERS_reg_11_39_inst : DLH_X1 port map( G => n11984, D => N3574, Q 
                           => NEXT_REGISTERS_11_39_port);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => N1341, CK => CLK, Q => 
                           n_1344, QN => n729_port);
   NEXT_REGISTERS_reg_11_38_inst : DLH_X1 port map( G => n11984, D => N3573, Q 
                           => NEXT_REGISTERS_11_38_port);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => N1340, CK => CLK, Q => 
                           n_1345, QN => n730_port);
   NEXT_REGISTERS_reg_11_37_inst : DLH_X1 port map( G => n11984, D => N3572, Q 
                           => NEXT_REGISTERS_11_37_port);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => N1339, CK => CLK, Q => 
                           n_1346, QN => n731_port);
   NEXT_REGISTERS_reg_11_36_inst : DLH_X1 port map( G => n11984, D => N3571, Q 
                           => NEXT_REGISTERS_11_36_port);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => N1338, CK => CLK, Q => 
                           n_1347, QN => n732_port);
   NEXT_REGISTERS_reg_11_35_inst : DLH_X1 port map( G => n11984, D => N3570, Q 
                           => NEXT_REGISTERS_11_35_port);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => N1337, CK => CLK, Q => 
                           n_1348, QN => n733_port);
   NEXT_REGISTERS_reg_11_34_inst : DLH_X1 port map( G => n11984, D => N3569, Q 
                           => NEXT_REGISTERS_11_34_port);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => N1336, CK => CLK, Q => 
                           n_1349, QN => n734_port);
   NEXT_REGISTERS_reg_11_33_inst : DLH_X1 port map( G => n11984, D => N3568, Q 
                           => NEXT_REGISTERS_11_33_port);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => N1335, CK => CLK, Q => 
                           n_1350, QN => n735_port);
   NEXT_REGISTERS_reg_11_32_inst : DLH_X1 port map( G => n11984, D => N3567, Q 
                           => NEXT_REGISTERS_11_32_port);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => N1334, CK => CLK, Q => 
                           n_1351, QN => n736_port);
   NEXT_REGISTERS_reg_11_31_inst : DLH_X1 port map( G => n11984, D => N3566, Q 
                           => NEXT_REGISTERS_11_31_port);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => N1333, CK => CLK, Q => 
                           n_1352, QN => n737_port);
   NEXT_REGISTERS_reg_11_30_inst : DLH_X1 port map( G => n11985, D => N3565, Q 
                           => NEXT_REGISTERS_11_30_port);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => N1332, CK => CLK, Q => 
                           n_1353, QN => n738_port);
   NEXT_REGISTERS_reg_11_29_inst : DLH_X1 port map( G => n11985, D => N3564, Q 
                           => NEXT_REGISTERS_11_29_port);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => N1331, CK => CLK, Q => 
                           n_1354, QN => n739_port);
   NEXT_REGISTERS_reg_11_28_inst : DLH_X1 port map( G => n11985, D => N3563, Q 
                           => NEXT_REGISTERS_11_28_port);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => N1330, CK => CLK, Q => 
                           n_1355, QN => n740_port);
   NEXT_REGISTERS_reg_11_27_inst : DLH_X1 port map( G => n11985, D => N3562, Q 
                           => NEXT_REGISTERS_11_27_port);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => N1329, CK => CLK, Q => 
                           n_1356, QN => n741_port);
   NEXT_REGISTERS_reg_11_26_inst : DLH_X1 port map( G => n11985, D => N3561, Q 
                           => NEXT_REGISTERS_11_26_port);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => N1328, CK => CLK, Q => 
                           n_1357, QN => n742_port);
   NEXT_REGISTERS_reg_11_25_inst : DLH_X1 port map( G => n11985, D => N3560, Q 
                           => NEXT_REGISTERS_11_25_port);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => N1327, CK => CLK, Q => 
                           n_1358, QN => n743_port);
   NEXT_REGISTERS_reg_11_24_inst : DLH_X1 port map( G => n11985, D => N3559, Q 
                           => NEXT_REGISTERS_11_24_port);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => N1326, CK => CLK, Q => 
                           n_1359, QN => n744_port);
   NEXT_REGISTERS_reg_11_23_inst : DLH_X1 port map( G => n11985, D => N3558, Q 
                           => NEXT_REGISTERS_11_23_port);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => N1325, CK => CLK, Q => 
                           n_1360, QN => n745_port);
   NEXT_REGISTERS_reg_11_22_inst : DLH_X1 port map( G => n11985, D => N3557, Q 
                           => NEXT_REGISTERS_11_22_port);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => N1324, CK => CLK, Q => 
                           n_1361, QN => n746_port);
   NEXT_REGISTERS_reg_11_21_inst : DLH_X1 port map( G => n11985, D => N3556, Q 
                           => NEXT_REGISTERS_11_21_port);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => N1323, CK => CLK, Q => 
                           n_1362, QN => n747_port);
   NEXT_REGISTERS_reg_11_20_inst : DLH_X1 port map( G => n11985, D => N3555, Q 
                           => NEXT_REGISTERS_11_20_port);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => N1322, CK => CLK, Q => 
                           n_1363, QN => n748_port);
   NEXT_REGISTERS_reg_11_19_inst : DLH_X1 port map( G => n11986, D => N3554, Q 
                           => NEXT_REGISTERS_11_19_port);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => N1321, CK => CLK, Q => 
                           n_1364, QN => n749_port);
   NEXT_REGISTERS_reg_11_18_inst : DLH_X1 port map( G => n11986, D => N3553, Q 
                           => NEXT_REGISTERS_11_18_port);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => N1320, CK => CLK, Q => 
                           n_1365, QN => n750_port);
   NEXT_REGISTERS_reg_11_17_inst : DLH_X1 port map( G => n11986, D => N3552, Q 
                           => NEXT_REGISTERS_11_17_port);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => N1319, CK => CLK, Q => 
                           n_1366, QN => n751_port);
   NEXT_REGISTERS_reg_11_16_inst : DLH_X1 port map( G => n11986, D => N3551, Q 
                           => NEXT_REGISTERS_11_16_port);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => N1318, CK => CLK, Q => 
                           n_1367, QN => n752_port);
   NEXT_REGISTERS_reg_11_15_inst : DLH_X1 port map( G => n11986, D => N3550, Q 
                           => NEXT_REGISTERS_11_15_port);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => N1317, CK => CLK, Q => 
                           n_1368, QN => n753_port);
   NEXT_REGISTERS_reg_11_14_inst : DLH_X1 port map( G => n11986, D => N3549, Q 
                           => NEXT_REGISTERS_11_14_port);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => N1316, CK => CLK, Q => 
                           n_1369, QN => n754_port);
   NEXT_REGISTERS_reg_11_13_inst : DLH_X1 port map( G => n11986, D => N3548, Q 
                           => NEXT_REGISTERS_11_13_port);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => N1315, CK => CLK, Q => 
                           n_1370, QN => n755_port);
   NEXT_REGISTERS_reg_11_12_inst : DLH_X1 port map( G => n11986, D => N3547, Q 
                           => NEXT_REGISTERS_11_12_port);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => N1314, CK => CLK, Q => 
                           n_1371, QN => n756_port);
   NEXT_REGISTERS_reg_11_11_inst : DLH_X1 port map( G => n11986, D => N3546, Q 
                           => NEXT_REGISTERS_11_11_port);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => N1313, CK => CLK, Q => 
                           n_1372, QN => n757_port);
   NEXT_REGISTERS_reg_11_10_inst : DLH_X1 port map( G => n11986, D => N3545, Q 
                           => NEXT_REGISTERS_11_10_port);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => N1312, CK => CLK, Q => 
                           n_1373, QN => n758_port);
   NEXT_REGISTERS_reg_11_9_inst : DLH_X1 port map( G => n11986, D => N3544, Q 
                           => NEXT_REGISTERS_11_9_port);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => N1311, CK => CLK, Q => 
                           n_1374, QN => n759_port);
   NEXT_REGISTERS_reg_11_8_inst : DLH_X1 port map( G => n11987, D => N3543, Q 
                           => NEXT_REGISTERS_11_8_port);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => N1310, CK => CLK, Q => 
                           n_1375, QN => n760_port);
   NEXT_REGISTERS_reg_11_7_inst : DLH_X1 port map( G => n11987, D => N3542, Q 
                           => NEXT_REGISTERS_11_7_port);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => N1309, CK => CLK, Q => 
                           n_1376, QN => n761_port);
   NEXT_REGISTERS_reg_11_6_inst : DLH_X1 port map( G => n11987, D => N3541, Q 
                           => NEXT_REGISTERS_11_6_port);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => N1308, CK => CLK, Q => 
                           n_1377, QN => n762_port);
   NEXT_REGISTERS_reg_11_5_inst : DLH_X1 port map( G => n11987, D => N3540, Q 
                           => NEXT_REGISTERS_11_5_port);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => N1307, CK => CLK, Q => 
                           n_1378, QN => n763_port);
   NEXT_REGISTERS_reg_11_4_inst : DLH_X1 port map( G => n11987, D => N3539, Q 
                           => NEXT_REGISTERS_11_4_port);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => N1306, CK => CLK, Q => 
                           n_1379, QN => n764_port);
   NEXT_REGISTERS_reg_11_3_inst : DLH_X1 port map( G => n11987, D => N3538, Q 
                           => NEXT_REGISTERS_11_3_port);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => N1305, CK => CLK, Q => 
                           n_1380, QN => n765_port);
   NEXT_REGISTERS_reg_11_2_inst : DLH_X1 port map( G => n11987, D => N3537, Q 
                           => NEXT_REGISTERS_11_2_port);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => N1304, CK => CLK, Q => 
                           n_1381, QN => n766_port);
   NEXT_REGISTERS_reg_11_1_inst : DLH_X1 port map( G => n11987, D => N3536, Q 
                           => NEXT_REGISTERS_11_1_port);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => N1303, CK => CLK, Q => 
                           n_1382, QN => n767_port);
   NEXT_REGISTERS_reg_11_0_inst : DLH_X1 port map( G => n11987, D => N3535, Q 
                           => NEXT_REGISTERS_11_0_port);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => N1302, CK => CLK, Q => 
                           n_1383, QN => n768_port);
   NEXT_REGISTERS_reg_12_63_inst : DLH_X1 port map( G => n11991, D => N3533, Q 
                           => NEXT_REGISTERS_12_63_port);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => N1301, CK => CLK, Q => 
                           n_1384, QN => n769_port);
   NEXT_REGISTERS_reg_12_62_inst : DLH_X1 port map( G => n11991, D => N3532, Q 
                           => NEXT_REGISTERS_12_62_port);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => N1300, CK => CLK, Q => 
                           n_1385, QN => n770_port);
   NEXT_REGISTERS_reg_12_61_inst : DLH_X1 port map( G => n11991, D => N3531, Q 
                           => NEXT_REGISTERS_12_61_port);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => N1299, CK => CLK, Q => 
                           n_1386, QN => n771_port);
   NEXT_REGISTERS_reg_12_60_inst : DLH_X1 port map( G => n11991, D => N3530, Q 
                           => NEXT_REGISTERS_12_60_port);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => N1298, CK => CLK, Q => 
                           n_1387, QN => n772_port);
   NEXT_REGISTERS_reg_12_59_inst : DLH_X1 port map( G => n11991, D => N3529, Q 
                           => NEXT_REGISTERS_12_59_port);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => N1297, CK => CLK, Q => 
                           n_1388, QN => n773_port);
   NEXT_REGISTERS_reg_12_58_inst : DLH_X1 port map( G => n11991, D => N3528, Q 
                           => NEXT_REGISTERS_12_58_port);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => N1296, CK => CLK, Q => 
                           n_1389, QN => n774_port);
   NEXT_REGISTERS_reg_12_57_inst : DLH_X1 port map( G => n11991, D => N3527, Q 
                           => NEXT_REGISTERS_12_57_port);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => N1295, CK => CLK, Q => 
                           n_1390, QN => n775_port);
   NEXT_REGISTERS_reg_12_56_inst : DLH_X1 port map( G => n11991, D => N3526, Q 
                           => NEXT_REGISTERS_12_56_port);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => N1294, CK => CLK, Q => 
                           n_1391, QN => n776_port);
   NEXT_REGISTERS_reg_12_55_inst : DLH_X1 port map( G => n11991, D => N3525, Q 
                           => NEXT_REGISTERS_12_55_port);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => N1293, CK => CLK, Q => 
                           n_1392, QN => n777_port);
   NEXT_REGISTERS_reg_12_54_inst : DLH_X1 port map( G => n11991, D => N3524, Q 
                           => NEXT_REGISTERS_12_54_port);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => N1292, CK => CLK, Q => 
                           n_1393, QN => n778_port);
   NEXT_REGISTERS_reg_12_53_inst : DLH_X1 port map( G => n11991, D => N3523, Q 
                           => NEXT_REGISTERS_12_53_port);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => N1291, CK => CLK, Q => 
                           n_1394, QN => n779_port);
   NEXT_REGISTERS_reg_12_52_inst : DLH_X1 port map( G => n11992, D => N3522, Q 
                           => NEXT_REGISTERS_12_52_port);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => N1290, CK => CLK, Q => 
                           n_1395, QN => n780_port);
   NEXT_REGISTERS_reg_12_51_inst : DLH_X1 port map( G => n11992, D => N3521, Q 
                           => NEXT_REGISTERS_12_51_port);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => N1289, CK => CLK, Q => 
                           n_1396, QN => n781_port);
   NEXT_REGISTERS_reg_12_50_inst : DLH_X1 port map( G => n11992, D => N3520, Q 
                           => NEXT_REGISTERS_12_50_port);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => N1288, CK => CLK, Q => 
                           n_1397, QN => n782_port);
   NEXT_REGISTERS_reg_12_49_inst : DLH_X1 port map( G => n11992, D => N3519, Q 
                           => NEXT_REGISTERS_12_49_port);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => N1287, CK => CLK, Q => 
                           n_1398, QN => n783_port);
   NEXT_REGISTERS_reg_12_48_inst : DLH_X1 port map( G => n11992, D => N3518, Q 
                           => NEXT_REGISTERS_12_48_port);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => N1286, CK => CLK, Q => 
                           n_1399, QN => n784_port);
   NEXT_REGISTERS_reg_12_47_inst : DLH_X1 port map( G => n11992, D => N3517, Q 
                           => NEXT_REGISTERS_12_47_port);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => N1285, CK => CLK, Q => 
                           n_1400, QN => n785_port);
   NEXT_REGISTERS_reg_12_46_inst : DLH_X1 port map( G => n11992, D => N3516, Q 
                           => NEXT_REGISTERS_12_46_port);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => N1284, CK => CLK, Q => 
                           n_1401, QN => n786_port);
   NEXT_REGISTERS_reg_12_45_inst : DLH_X1 port map( G => n11992, D => N3515, Q 
                           => NEXT_REGISTERS_12_45_port);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => N1283, CK => CLK, Q => 
                           n_1402, QN => n787_port);
   NEXT_REGISTERS_reg_12_44_inst : DLH_X1 port map( G => n11992, D => N3514, Q 
                           => NEXT_REGISTERS_12_44_port);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => N1282, CK => CLK, Q => 
                           n_1403, QN => n788_port);
   NEXT_REGISTERS_reg_12_43_inst : DLH_X1 port map( G => n11992, D => N3513, Q 
                           => NEXT_REGISTERS_12_43_port);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => N1281, CK => CLK, Q => 
                           n_1404, QN => n789_port);
   NEXT_REGISTERS_reg_12_42_inst : DLH_X1 port map( G => n11992, D => N3512, Q 
                           => NEXT_REGISTERS_12_42_port);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => N1280, CK => CLK, Q => 
                           n_1405, QN => n790_port);
   NEXT_REGISTERS_reg_12_41_inst : DLH_X1 port map( G => n11993, D => N3511, Q 
                           => NEXT_REGISTERS_12_41_port);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => N1279, CK => CLK, Q => 
                           n_1406, QN => n791_port);
   NEXT_REGISTERS_reg_12_40_inst : DLH_X1 port map( G => n11993, D => N3510, Q 
                           => NEXT_REGISTERS_12_40_port);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => N1278, CK => CLK, Q => 
                           n_1407, QN => n792_port);
   NEXT_REGISTERS_reg_12_39_inst : DLH_X1 port map( G => n11993, D => N3509, Q 
                           => NEXT_REGISTERS_12_39_port);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => N1277, CK => CLK, Q => 
                           n_1408, QN => n793_port);
   NEXT_REGISTERS_reg_12_38_inst : DLH_X1 port map( G => n11993, D => N3508, Q 
                           => NEXT_REGISTERS_12_38_port);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => N1276, CK => CLK, Q => 
                           n_1409, QN => n794_port);
   NEXT_REGISTERS_reg_12_37_inst : DLH_X1 port map( G => n11993, D => N3507, Q 
                           => NEXT_REGISTERS_12_37_port);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => N1275, CK => CLK, Q => 
                           n_1410, QN => n795_port);
   NEXT_REGISTERS_reg_12_36_inst : DLH_X1 port map( G => n11993, D => N3506, Q 
                           => NEXT_REGISTERS_12_36_port);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => N1274, CK => CLK, Q => 
                           n_1411, QN => n796_port);
   NEXT_REGISTERS_reg_12_35_inst : DLH_X1 port map( G => n11993, D => N3505, Q 
                           => NEXT_REGISTERS_12_35_port);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => N1273, CK => CLK, Q => 
                           n_1412, QN => n797_port);
   NEXT_REGISTERS_reg_12_34_inst : DLH_X1 port map( G => n11993, D => N3504, Q 
                           => NEXT_REGISTERS_12_34_port);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => N1272, CK => CLK, Q => 
                           n_1413, QN => n798_port);
   NEXT_REGISTERS_reg_12_33_inst : DLH_X1 port map( G => n11993, D => N3503, Q 
                           => NEXT_REGISTERS_12_33_port);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => N1271, CK => CLK, Q => 
                           n_1414, QN => n799_port);
   NEXT_REGISTERS_reg_12_32_inst : DLH_X1 port map( G => n11993, D => N3502, Q 
                           => NEXT_REGISTERS_12_32_port);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => N1270, CK => CLK, Q => 
                           n_1415, QN => n800_port);
   NEXT_REGISTERS_reg_12_31_inst : DLH_X1 port map( G => n11993, D => N3501, Q 
                           => NEXT_REGISTERS_12_31_port);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => N1269, CK => CLK, Q => 
                           n_1416, QN => n801_port);
   NEXT_REGISTERS_reg_12_30_inst : DLH_X1 port map( G => n11994, D => N3500, Q 
                           => NEXT_REGISTERS_12_30_port);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => N1268, CK => CLK, Q => 
                           n_1417, QN => n802_port);
   NEXT_REGISTERS_reg_12_29_inst : DLH_X1 port map( G => n11994, D => N3499, Q 
                           => NEXT_REGISTERS_12_29_port);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => N1267, CK => CLK, Q => 
                           n_1418, QN => n803_port);
   NEXT_REGISTERS_reg_12_28_inst : DLH_X1 port map( G => n11994, D => N3498, Q 
                           => NEXT_REGISTERS_12_28_port);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => N1266, CK => CLK, Q => 
                           n_1419, QN => n804_port);
   NEXT_REGISTERS_reg_12_27_inst : DLH_X1 port map( G => n11994, D => N3497, Q 
                           => NEXT_REGISTERS_12_27_port);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => N1265, CK => CLK, Q => 
                           n_1420, QN => n805_port);
   NEXT_REGISTERS_reg_12_26_inst : DLH_X1 port map( G => n11994, D => N3496, Q 
                           => NEXT_REGISTERS_12_26_port);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => N1264, CK => CLK, Q => 
                           n_1421, QN => n806_port);
   NEXT_REGISTERS_reg_12_25_inst : DLH_X1 port map( G => n11994, D => N3495, Q 
                           => NEXT_REGISTERS_12_25_port);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => N1263, CK => CLK, Q => 
                           n_1422, QN => n807_port);
   NEXT_REGISTERS_reg_12_24_inst : DLH_X1 port map( G => n11994, D => N3494, Q 
                           => NEXT_REGISTERS_12_24_port);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => N1262, CK => CLK, Q => 
                           n_1423, QN => n808_port);
   NEXT_REGISTERS_reg_12_23_inst : DLH_X1 port map( G => n11994, D => N3493, Q 
                           => NEXT_REGISTERS_12_23_port);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => N1261, CK => CLK, Q => 
                           n_1424, QN => n809_port);
   NEXT_REGISTERS_reg_12_22_inst : DLH_X1 port map( G => n11994, D => N3492, Q 
                           => NEXT_REGISTERS_12_22_port);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => N1260, CK => CLK, Q => 
                           n_1425, QN => n810_port);
   NEXT_REGISTERS_reg_12_21_inst : DLH_X1 port map( G => n11994, D => N3491, Q 
                           => NEXT_REGISTERS_12_21_port);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => N1259, CK => CLK, Q => 
                           n_1426, QN => n811_port);
   NEXT_REGISTERS_reg_12_20_inst : DLH_X1 port map( G => n11994, D => N3490, Q 
                           => NEXT_REGISTERS_12_20_port);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => N1258, CK => CLK, Q => 
                           n_1427, QN => n812_port);
   NEXT_REGISTERS_reg_12_19_inst : DLH_X1 port map( G => n11995, D => N3489, Q 
                           => NEXT_REGISTERS_12_19_port);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => N1257, CK => CLK, Q => 
                           n_1428, QN => n813_port);
   NEXT_REGISTERS_reg_12_18_inst : DLH_X1 port map( G => n11995, D => N3488, Q 
                           => NEXT_REGISTERS_12_18_port);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => N1256, CK => CLK, Q => 
                           n_1429, QN => n814_port);
   NEXT_REGISTERS_reg_12_17_inst : DLH_X1 port map( G => n11995, D => N3487, Q 
                           => NEXT_REGISTERS_12_17_port);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => N1255, CK => CLK, Q => 
                           n_1430, QN => n815_port);
   NEXT_REGISTERS_reg_12_16_inst : DLH_X1 port map( G => n11995, D => N3486, Q 
                           => NEXT_REGISTERS_12_16_port);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => N1254, CK => CLK, Q => 
                           n_1431, QN => n816_port);
   NEXT_REGISTERS_reg_12_15_inst : DLH_X1 port map( G => n11995, D => N3485, Q 
                           => NEXT_REGISTERS_12_15_port);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => N1253, CK => CLK, Q => 
                           n_1432, QN => n817_port);
   NEXT_REGISTERS_reg_12_14_inst : DLH_X1 port map( G => n11995, D => N3484, Q 
                           => NEXT_REGISTERS_12_14_port);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => N1252, CK => CLK, Q => 
                           n_1433, QN => n818_port);
   NEXT_REGISTERS_reg_12_13_inst : DLH_X1 port map( G => n11995, D => N3483, Q 
                           => NEXT_REGISTERS_12_13_port);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => N1251, CK => CLK, Q => 
                           n_1434, QN => n819_port);
   NEXT_REGISTERS_reg_12_12_inst : DLH_X1 port map( G => n11995, D => N3482, Q 
                           => NEXT_REGISTERS_12_12_port);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => N1250, CK => CLK, Q => 
                           n_1435, QN => n820_port);
   NEXT_REGISTERS_reg_12_11_inst : DLH_X1 port map( G => n11995, D => N3481, Q 
                           => NEXT_REGISTERS_12_11_port);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => N1249, CK => CLK, Q => 
                           n_1436, QN => n821_port);
   NEXT_REGISTERS_reg_12_10_inst : DLH_X1 port map( G => n11995, D => N3480, Q 
                           => NEXT_REGISTERS_12_10_port);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => N1248, CK => CLK, Q => 
                           n_1437, QN => n822_port);
   NEXT_REGISTERS_reg_12_9_inst : DLH_X1 port map( G => n11995, D => N3479, Q 
                           => NEXT_REGISTERS_12_9_port);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => N1247, CK => CLK, Q => 
                           n_1438, QN => n823_port);
   NEXT_REGISTERS_reg_12_8_inst : DLH_X1 port map( G => n11996, D => N3478, Q 
                           => NEXT_REGISTERS_12_8_port);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => N1246, CK => CLK, Q => 
                           n_1439, QN => n824_port);
   NEXT_REGISTERS_reg_12_7_inst : DLH_X1 port map( G => n11996, D => N3477, Q 
                           => NEXT_REGISTERS_12_7_port);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => N1245, CK => CLK, Q => 
                           n_1440, QN => n825_port);
   NEXT_REGISTERS_reg_12_6_inst : DLH_X1 port map( G => n11996, D => N3476, Q 
                           => NEXT_REGISTERS_12_6_port);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => N1244, CK => CLK, Q => 
                           n_1441, QN => n826_port);
   NEXT_REGISTERS_reg_12_5_inst : DLH_X1 port map( G => n11996, D => N3475, Q 
                           => NEXT_REGISTERS_12_5_port);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => N1243, CK => CLK, Q => 
                           n_1442, QN => n827_port);
   NEXT_REGISTERS_reg_12_4_inst : DLH_X1 port map( G => n11996, D => N3474, Q 
                           => NEXT_REGISTERS_12_4_port);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => N1242, CK => CLK, Q => 
                           n_1443, QN => n828_port);
   NEXT_REGISTERS_reg_12_3_inst : DLH_X1 port map( G => n11996, D => N3473, Q 
                           => NEXT_REGISTERS_12_3_port);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => N1241, CK => CLK, Q => 
                           n_1444, QN => n829_port);
   NEXT_REGISTERS_reg_12_2_inst : DLH_X1 port map( G => n11996, D => N3472, Q 
                           => NEXT_REGISTERS_12_2_port);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => N1240, CK => CLK, Q => 
                           n_1445, QN => n830_port);
   NEXT_REGISTERS_reg_12_1_inst : DLH_X1 port map( G => n11996, D => N3471, Q 
                           => NEXT_REGISTERS_12_1_port);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => N1239, CK => CLK, Q => 
                           n_1446, QN => n831_port);
   NEXT_REGISTERS_reg_12_0_inst : DLH_X1 port map( G => n11996, D => N3470, Q 
                           => NEXT_REGISTERS_12_0_port);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => N1238, CK => CLK, Q => 
                           n_1447, QN => n832_port);
   NEXT_REGISTERS_reg_13_63_inst : DLH_X1 port map( G => n12000, D => N3468, Q 
                           => NEXT_REGISTERS_13_63_port);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => N1237, CK => CLK, Q => 
                           n10093, QN => n833_port);
   NEXT_REGISTERS_reg_13_62_inst : DLH_X1 port map( G => n12000, D => N3467, Q 
                           => NEXT_REGISTERS_13_62_port);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => N1236, CK => CLK, Q => 
                           n10091, QN => n834_port);
   NEXT_REGISTERS_reg_13_61_inst : DLH_X1 port map( G => n12000, D => N3466, Q 
                           => NEXT_REGISTERS_13_61_port);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => N1235, CK => CLK, Q => 
                           n10089, QN => n835_port);
   NEXT_REGISTERS_reg_13_60_inst : DLH_X1 port map( G => n12000, D => N3465, Q 
                           => NEXT_REGISTERS_13_60_port);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => N1234, CK => CLK, Q => 
                           n10087, QN => n836_port);
   NEXT_REGISTERS_reg_13_59_inst : DLH_X1 port map( G => n12000, D => N3464, Q 
                           => NEXT_REGISTERS_13_59_port);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => N1233, CK => CLK, Q => 
                           n10085, QN => n837_port);
   NEXT_REGISTERS_reg_13_58_inst : DLH_X1 port map( G => n12000, D => N3463, Q 
                           => NEXT_REGISTERS_13_58_port);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => N1232, CK => CLK, Q => 
                           n10083, QN => n838_port);
   NEXT_REGISTERS_reg_13_57_inst : DLH_X1 port map( G => n12000, D => N3462, Q 
                           => NEXT_REGISTERS_13_57_port);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => N1231, CK => CLK, Q => 
                           n10081, QN => n839_port);
   NEXT_REGISTERS_reg_13_56_inst : DLH_X1 port map( G => n12000, D => N3461, Q 
                           => NEXT_REGISTERS_13_56_port);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => N1230, CK => CLK, Q => 
                           n10079, QN => n840_port);
   NEXT_REGISTERS_reg_13_55_inst : DLH_X1 port map( G => n12000, D => N3460, Q 
                           => NEXT_REGISTERS_13_55_port);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => N1229, CK => CLK, Q => 
                           n10077, QN => n841_port);
   NEXT_REGISTERS_reg_13_54_inst : DLH_X1 port map( G => n12000, D => N3459, Q 
                           => NEXT_REGISTERS_13_54_port);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => N1228, CK => CLK, Q => 
                           n10075, QN => n842_port);
   NEXT_REGISTERS_reg_13_53_inst : DLH_X1 port map( G => n12000, D => N3458, Q 
                           => NEXT_REGISTERS_13_53_port);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => N1227, CK => CLK, Q => 
                           n10073, QN => n843_port);
   NEXT_REGISTERS_reg_13_52_inst : DLH_X1 port map( G => n12001, D => N3457, Q 
                           => NEXT_REGISTERS_13_52_port);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => N1226, CK => CLK, Q => 
                           n10071, QN => n844_port);
   NEXT_REGISTERS_reg_13_51_inst : DLH_X1 port map( G => n12001, D => N3456, Q 
                           => NEXT_REGISTERS_13_51_port);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => N1225, CK => CLK, Q => 
                           n10069, QN => n845_port);
   NEXT_REGISTERS_reg_13_50_inst : DLH_X1 port map( G => n12001, D => N3455, Q 
                           => NEXT_REGISTERS_13_50_port);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => N1224, CK => CLK, Q => 
                           n10067, QN => n846_port);
   NEXT_REGISTERS_reg_13_49_inst : DLH_X1 port map( G => n12001, D => N3454, Q 
                           => NEXT_REGISTERS_13_49_port);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => N1223, CK => CLK, Q => 
                           n10065, QN => n847_port);
   NEXT_REGISTERS_reg_13_48_inst : DLH_X1 port map( G => n12001, D => N3453, Q 
                           => NEXT_REGISTERS_13_48_port);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => N1222, CK => CLK, Q => 
                           n10063, QN => n848_port);
   NEXT_REGISTERS_reg_13_47_inst : DLH_X1 port map( G => n12001, D => N3452, Q 
                           => NEXT_REGISTERS_13_47_port);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => N1221, CK => CLK, Q => 
                           n10061, QN => n849_port);
   NEXT_REGISTERS_reg_13_46_inst : DLH_X1 port map( G => n12001, D => N3451, Q 
                           => NEXT_REGISTERS_13_46_port);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => N1220, CK => CLK, Q => 
                           n10059, QN => n850_port);
   NEXT_REGISTERS_reg_13_45_inst : DLH_X1 port map( G => n12001, D => N3450, Q 
                           => NEXT_REGISTERS_13_45_port);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => N1219, CK => CLK, Q => 
                           n10057, QN => n851_port);
   NEXT_REGISTERS_reg_13_44_inst : DLH_X1 port map( G => n12001, D => N3449, Q 
                           => NEXT_REGISTERS_13_44_port);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => N1218, CK => CLK, Q => 
                           n10055, QN => n852_port);
   NEXT_REGISTERS_reg_13_43_inst : DLH_X1 port map( G => n12001, D => N3448, Q 
                           => NEXT_REGISTERS_13_43_port);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => N1217, CK => CLK, Q => 
                           n10053, QN => n853_port);
   NEXT_REGISTERS_reg_13_42_inst : DLH_X1 port map( G => n12001, D => N3447, Q 
                           => NEXT_REGISTERS_13_42_port);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => N1216, CK => CLK, Q => 
                           n10051, QN => n854_port);
   NEXT_REGISTERS_reg_13_41_inst : DLH_X1 port map( G => n12002, D => N3446, Q 
                           => NEXT_REGISTERS_13_41_port);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => N1215, CK => CLK, Q => 
                           n10049, QN => n855_port);
   NEXT_REGISTERS_reg_13_40_inst : DLH_X1 port map( G => n12002, D => N3445, Q 
                           => NEXT_REGISTERS_13_40_port);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => N1214, CK => CLK, Q => 
                           n10047, QN => n856_port);
   NEXT_REGISTERS_reg_13_39_inst : DLH_X1 port map( G => n12002, D => N3444, Q 
                           => NEXT_REGISTERS_13_39_port);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => N1213, CK => CLK, Q => 
                           n10045, QN => n857_port);
   NEXT_REGISTERS_reg_13_38_inst : DLH_X1 port map( G => n12002, D => N3443, Q 
                           => NEXT_REGISTERS_13_38_port);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => N1212, CK => CLK, Q => 
                           n10043, QN => n858_port);
   NEXT_REGISTERS_reg_13_37_inst : DLH_X1 port map( G => n12002, D => N3442, Q 
                           => NEXT_REGISTERS_13_37_port);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => N1211, CK => CLK, Q => 
                           n10041, QN => n859_port);
   NEXT_REGISTERS_reg_13_36_inst : DLH_X1 port map( G => n12002, D => N3441, Q 
                           => NEXT_REGISTERS_13_36_port);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => N1210, CK => CLK, Q => 
                           n10039, QN => n860_port);
   NEXT_REGISTERS_reg_13_35_inst : DLH_X1 port map( G => n12002, D => N3440, Q 
                           => NEXT_REGISTERS_13_35_port);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => N1209, CK => CLK, Q => 
                           n10037, QN => n861_port);
   NEXT_REGISTERS_reg_13_34_inst : DLH_X1 port map( G => n12002, D => N3439, Q 
                           => NEXT_REGISTERS_13_34_port);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => N1208, CK => CLK, Q => 
                           n10035, QN => n862_port);
   NEXT_REGISTERS_reg_13_33_inst : DLH_X1 port map( G => n12002, D => N3438, Q 
                           => NEXT_REGISTERS_13_33_port);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => N1207, CK => CLK, Q => 
                           n10033, QN => n863_port);
   NEXT_REGISTERS_reg_13_32_inst : DLH_X1 port map( G => n12002, D => N3437, Q 
                           => NEXT_REGISTERS_13_32_port);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => N1206, CK => CLK, Q => 
                           n10031, QN => n864_port);
   NEXT_REGISTERS_reg_13_31_inst : DLH_X1 port map( G => n12002, D => N3436, Q 
                           => NEXT_REGISTERS_13_31_port);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => N1205, CK => CLK, Q => 
                           n10029, QN => n865_port);
   NEXT_REGISTERS_reg_13_30_inst : DLH_X1 port map( G => n12003, D => N3435, Q 
                           => NEXT_REGISTERS_13_30_port);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => N1204, CK => CLK, Q => 
                           n10027, QN => n866_port);
   NEXT_REGISTERS_reg_13_29_inst : DLH_X1 port map( G => n12003, D => N3434, Q 
                           => NEXT_REGISTERS_13_29_port);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => N1203, CK => CLK, Q => 
                           n10025, QN => n867_port);
   NEXT_REGISTERS_reg_13_28_inst : DLH_X1 port map( G => n12003, D => N3433, Q 
                           => NEXT_REGISTERS_13_28_port);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => N1202, CK => CLK, Q => 
                           n10023, QN => n868_port);
   NEXT_REGISTERS_reg_13_27_inst : DLH_X1 port map( G => n12003, D => N3432, Q 
                           => NEXT_REGISTERS_13_27_port);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => N1201, CK => CLK, Q => 
                           n10021, QN => n869_port);
   NEXT_REGISTERS_reg_13_26_inst : DLH_X1 port map( G => n12003, D => N3431, Q 
                           => NEXT_REGISTERS_13_26_port);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => N1200, CK => CLK, Q => 
                           n10019, QN => n870_port);
   NEXT_REGISTERS_reg_13_25_inst : DLH_X1 port map( G => n12003, D => N3430, Q 
                           => NEXT_REGISTERS_13_25_port);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => N1199, CK => CLK, Q => 
                           n10017, QN => n871_port);
   NEXT_REGISTERS_reg_13_24_inst : DLH_X1 port map( G => n12003, D => N3429, Q 
                           => NEXT_REGISTERS_13_24_port);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => N1198, CK => CLK, Q => 
                           n10015, QN => n872_port);
   NEXT_REGISTERS_reg_13_23_inst : DLH_X1 port map( G => n12003, D => N3428, Q 
                           => NEXT_REGISTERS_13_23_port);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => N1197, CK => CLK, Q => 
                           n10013, QN => n873_port);
   NEXT_REGISTERS_reg_13_22_inst : DLH_X1 port map( G => n12003, D => N3427, Q 
                           => NEXT_REGISTERS_13_22_port);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => N1196, CK => CLK, Q => 
                           n10011, QN => n874_port);
   NEXT_REGISTERS_reg_13_21_inst : DLH_X1 port map( G => n12003, D => N3426, Q 
                           => NEXT_REGISTERS_13_21_port);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => N1195, CK => CLK, Q => 
                           n10009, QN => n875_port);
   NEXT_REGISTERS_reg_13_20_inst : DLH_X1 port map( G => n12003, D => N3425, Q 
                           => NEXT_REGISTERS_13_20_port);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => N1194, CK => CLK, Q => 
                           n10007, QN => n876_port);
   NEXT_REGISTERS_reg_13_19_inst : DLH_X1 port map( G => n12004, D => N3424, Q 
                           => NEXT_REGISTERS_13_19_port);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => N1193, CK => CLK, Q => 
                           n10005, QN => n877_port);
   NEXT_REGISTERS_reg_13_18_inst : DLH_X1 port map( G => n12004, D => N3423, Q 
                           => NEXT_REGISTERS_13_18_port);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => N1192, CK => CLK, Q => 
                           n10003, QN => n878_port);
   NEXT_REGISTERS_reg_13_17_inst : DLH_X1 port map( G => n12004, D => N3422, Q 
                           => NEXT_REGISTERS_13_17_port);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => N1191, CK => CLK, Q => 
                           n10001, QN => n879_port);
   NEXT_REGISTERS_reg_13_16_inst : DLH_X1 port map( G => n12004, D => N3421, Q 
                           => NEXT_REGISTERS_13_16_port);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => N1190, CK => CLK, Q => 
                           n9999, QN => n880_port);
   NEXT_REGISTERS_reg_13_15_inst : DLH_X1 port map( G => n12004, D => N3420, Q 
                           => NEXT_REGISTERS_13_15_port);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => N1189, CK => CLK, Q => 
                           n9997, QN => n881_port);
   NEXT_REGISTERS_reg_13_14_inst : DLH_X1 port map( G => n12004, D => N3419, Q 
                           => NEXT_REGISTERS_13_14_port);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => N1188, CK => CLK, Q => 
                           n9995, QN => n882_port);
   NEXT_REGISTERS_reg_13_13_inst : DLH_X1 port map( G => n12004, D => N3418, Q 
                           => NEXT_REGISTERS_13_13_port);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => N1187, CK => CLK, Q => 
                           n9993, QN => n883_port);
   NEXT_REGISTERS_reg_13_12_inst : DLH_X1 port map( G => n12004, D => N3417, Q 
                           => NEXT_REGISTERS_13_12_port);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => N1186, CK => CLK, Q => 
                           n9991, QN => n884_port);
   NEXT_REGISTERS_reg_13_11_inst : DLH_X1 port map( G => n12004, D => N3416, Q 
                           => NEXT_REGISTERS_13_11_port);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => N1185, CK => CLK, Q => 
                           n9989, QN => n885_port);
   NEXT_REGISTERS_reg_13_10_inst : DLH_X1 port map( G => n12004, D => N3415, Q 
                           => NEXT_REGISTERS_13_10_port);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => N1184, CK => CLK, Q => 
                           n9987, QN => n886_port);
   NEXT_REGISTERS_reg_13_9_inst : DLH_X1 port map( G => n12004, D => N3414, Q 
                           => NEXT_REGISTERS_13_9_port);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => N1183, CK => CLK, Q => n9985
                           , QN => n887_port);
   NEXT_REGISTERS_reg_13_8_inst : DLH_X1 port map( G => n12005, D => N3413, Q 
                           => NEXT_REGISTERS_13_8_port);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => N1182, CK => CLK, Q => n9983
                           , QN => n888_port);
   NEXT_REGISTERS_reg_13_7_inst : DLH_X1 port map( G => n12005, D => N3412, Q 
                           => NEXT_REGISTERS_13_7_port);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => N1181, CK => CLK, Q => n9981
                           , QN => n889_port);
   NEXT_REGISTERS_reg_13_6_inst : DLH_X1 port map( G => n12005, D => N3411, Q 
                           => NEXT_REGISTERS_13_6_port);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => N1180, CK => CLK, Q => n9979
                           , QN => n890_port);
   NEXT_REGISTERS_reg_13_5_inst : DLH_X1 port map( G => n12005, D => N3410, Q 
                           => NEXT_REGISTERS_13_5_port);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => N1179, CK => CLK, Q => n9977
                           , QN => n891_port);
   NEXT_REGISTERS_reg_13_4_inst : DLH_X1 port map( G => n12005, D => N3409, Q 
                           => NEXT_REGISTERS_13_4_port);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => N1178, CK => CLK, Q => n9975
                           , QN => n892_port);
   NEXT_REGISTERS_reg_13_3_inst : DLH_X1 port map( G => n12005, D => N3408, Q 
                           => NEXT_REGISTERS_13_3_port);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => N1177, CK => CLK, Q => n9973
                           , QN => n893_port);
   NEXT_REGISTERS_reg_13_2_inst : DLH_X1 port map( G => n12005, D => N3407, Q 
                           => NEXT_REGISTERS_13_2_port);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => N1176, CK => CLK, Q => n9971
                           , QN => n894_port);
   NEXT_REGISTERS_reg_13_1_inst : DLH_X1 port map( G => n12005, D => N3406, Q 
                           => NEXT_REGISTERS_13_1_port);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => N1175, CK => CLK, Q => n9969
                           , QN => n895_port);
   NEXT_REGISTERS_reg_13_0_inst : DLH_X1 port map( G => n12005, D => N3405, Q 
                           => NEXT_REGISTERS_13_0_port);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => N1174, CK => CLK, Q => n9967
                           , QN => n896_port);
   NEXT_REGISTERS_reg_14_63_inst : DLH_X1 port map( G => n12009, D => N3403, Q 
                           => NEXT_REGISTERS_14_63_port);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => N1173, CK => CLK, Q => 
                           n_1448, QN => n897_port);
   NEXT_REGISTERS_reg_14_62_inst : DLH_X1 port map( G => n12009, D => N3402, Q 
                           => NEXT_REGISTERS_14_62_port);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => N1172, CK => CLK, Q => 
                           n_1449, QN => n898_port);
   NEXT_REGISTERS_reg_14_61_inst : DLH_X1 port map( G => n12009, D => N3401, Q 
                           => NEXT_REGISTERS_14_61_port);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => N1171, CK => CLK, Q => 
                           n_1450, QN => n899_port);
   NEXT_REGISTERS_reg_14_60_inst : DLH_X1 port map( G => n12009, D => N3400, Q 
                           => NEXT_REGISTERS_14_60_port);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => N1170, CK => CLK, Q => 
                           n_1451, QN => n900_port);
   NEXT_REGISTERS_reg_14_59_inst : DLH_X1 port map( G => n12009, D => N3399, Q 
                           => NEXT_REGISTERS_14_59_port);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => N1169, CK => CLK, Q => 
                           n_1452, QN => n901_port);
   NEXT_REGISTERS_reg_14_58_inst : DLH_X1 port map( G => n12009, D => N3398, Q 
                           => NEXT_REGISTERS_14_58_port);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => N1168, CK => CLK, Q => 
                           n_1453, QN => n902_port);
   NEXT_REGISTERS_reg_14_57_inst : DLH_X1 port map( G => n12009, D => N3397, Q 
                           => NEXT_REGISTERS_14_57_port);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => N1167, CK => CLK, Q => 
                           n_1454, QN => n903_port);
   NEXT_REGISTERS_reg_14_56_inst : DLH_X1 port map( G => n12009, D => N3396, Q 
                           => NEXT_REGISTERS_14_56_port);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => N1166, CK => CLK, Q => 
                           n_1455, QN => n904_port);
   NEXT_REGISTERS_reg_14_55_inst : DLH_X1 port map( G => n12009, D => N3395, Q 
                           => NEXT_REGISTERS_14_55_port);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => N1165, CK => CLK, Q => 
                           n_1456, QN => n905_port);
   NEXT_REGISTERS_reg_14_54_inst : DLH_X1 port map( G => n12009, D => N3394, Q 
                           => NEXT_REGISTERS_14_54_port);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => N1164, CK => CLK, Q => 
                           n_1457, QN => n906_port);
   NEXT_REGISTERS_reg_14_53_inst : DLH_X1 port map( G => n12009, D => N3393, Q 
                           => NEXT_REGISTERS_14_53_port);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => N1163, CK => CLK, Q => 
                           n_1458, QN => n907_port);
   NEXT_REGISTERS_reg_14_52_inst : DLH_X1 port map( G => n12010, D => N3392, Q 
                           => NEXT_REGISTERS_14_52_port);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => N1162, CK => CLK, Q => 
                           n_1459, QN => n908_port);
   NEXT_REGISTERS_reg_14_51_inst : DLH_X1 port map( G => n12010, D => N3391, Q 
                           => NEXT_REGISTERS_14_51_port);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => N1161, CK => CLK, Q => 
                           n_1460, QN => n909_port);
   NEXT_REGISTERS_reg_14_50_inst : DLH_X1 port map( G => n12010, D => N3390, Q 
                           => NEXT_REGISTERS_14_50_port);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => N1160, CK => CLK, Q => 
                           n_1461, QN => n910_port);
   NEXT_REGISTERS_reg_14_49_inst : DLH_X1 port map( G => n12010, D => N3389, Q 
                           => NEXT_REGISTERS_14_49_port);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => N1159, CK => CLK, Q => 
                           n_1462, QN => n911_port);
   NEXT_REGISTERS_reg_14_48_inst : DLH_X1 port map( G => n12010, D => N3388, Q 
                           => NEXT_REGISTERS_14_48_port);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => N1158, CK => CLK, Q => 
                           n_1463, QN => n912_port);
   NEXT_REGISTERS_reg_14_47_inst : DLH_X1 port map( G => n12010, D => N3387, Q 
                           => NEXT_REGISTERS_14_47_port);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => N1157, CK => CLK, Q => 
                           n_1464, QN => n913_port);
   NEXT_REGISTERS_reg_14_46_inst : DLH_X1 port map( G => n12010, D => N3386, Q 
                           => NEXT_REGISTERS_14_46_port);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => N1156, CK => CLK, Q => 
                           n_1465, QN => n914_port);
   NEXT_REGISTERS_reg_14_45_inst : DLH_X1 port map( G => n12010, D => N3385, Q 
                           => NEXT_REGISTERS_14_45_port);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => N1155, CK => CLK, Q => 
                           n_1466, QN => n915_port);
   NEXT_REGISTERS_reg_14_44_inst : DLH_X1 port map( G => n12010, D => N3384, Q 
                           => NEXT_REGISTERS_14_44_port);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => N1154, CK => CLK, Q => 
                           n_1467, QN => n916_port);
   NEXT_REGISTERS_reg_14_43_inst : DLH_X1 port map( G => n12010, D => N3383, Q 
                           => NEXT_REGISTERS_14_43_port);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => N1153, CK => CLK, Q => 
                           n_1468, QN => n917_port);
   NEXT_REGISTERS_reg_14_42_inst : DLH_X1 port map( G => n12010, D => N3382, Q 
                           => NEXT_REGISTERS_14_42_port);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => N1152, CK => CLK, Q => 
                           n_1469, QN => n918_port);
   NEXT_REGISTERS_reg_14_41_inst : DLH_X1 port map( G => n12011, D => N3381, Q 
                           => NEXT_REGISTERS_14_41_port);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => N1151, CK => CLK, Q => 
                           n_1470, QN => n919_port);
   NEXT_REGISTERS_reg_14_40_inst : DLH_X1 port map( G => n12011, D => N3380, Q 
                           => NEXT_REGISTERS_14_40_port);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => N1150, CK => CLK, Q => 
                           n_1471, QN => n920_port);
   NEXT_REGISTERS_reg_14_39_inst : DLH_X1 port map( G => n12011, D => N3379, Q 
                           => NEXT_REGISTERS_14_39_port);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => N1149, CK => CLK, Q => 
                           n_1472, QN => n921_port);
   NEXT_REGISTERS_reg_14_38_inst : DLH_X1 port map( G => n12011, D => N3378, Q 
                           => NEXT_REGISTERS_14_38_port);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => N1148, CK => CLK, Q => 
                           n_1473, QN => n922_port);
   NEXT_REGISTERS_reg_14_37_inst : DLH_X1 port map( G => n12011, D => N3377, Q 
                           => NEXT_REGISTERS_14_37_port);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => N1147, CK => CLK, Q => 
                           n_1474, QN => n923_port);
   NEXT_REGISTERS_reg_14_36_inst : DLH_X1 port map( G => n12011, D => N3376, Q 
                           => NEXT_REGISTERS_14_36_port);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => N1146, CK => CLK, Q => 
                           n_1475, QN => n924_port);
   NEXT_REGISTERS_reg_14_35_inst : DLH_X1 port map( G => n12011, D => N3375, Q 
                           => NEXT_REGISTERS_14_35_port);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => N1145, CK => CLK, Q => 
                           n_1476, QN => n925_port);
   NEXT_REGISTERS_reg_14_34_inst : DLH_X1 port map( G => n12011, D => N3374, Q 
                           => NEXT_REGISTERS_14_34_port);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => N1144, CK => CLK, Q => 
                           n_1477, QN => n926_port);
   NEXT_REGISTERS_reg_14_33_inst : DLH_X1 port map( G => n12011, D => N3373, Q 
                           => NEXT_REGISTERS_14_33_port);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => N1143, CK => CLK, Q => 
                           n_1478, QN => n927_port);
   NEXT_REGISTERS_reg_14_32_inst : DLH_X1 port map( G => n12011, D => N3372, Q 
                           => NEXT_REGISTERS_14_32_port);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => N1142, CK => CLK, Q => 
                           n_1479, QN => n928_port);
   NEXT_REGISTERS_reg_14_31_inst : DLH_X1 port map( G => n12011, D => N3371, Q 
                           => NEXT_REGISTERS_14_31_port);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => N1141, CK => CLK, Q => 
                           n_1480, QN => n929_port);
   NEXT_REGISTERS_reg_14_30_inst : DLH_X1 port map( G => n12012, D => N3370, Q 
                           => NEXT_REGISTERS_14_30_port);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => N1140, CK => CLK, Q => 
                           n_1481, QN => n930_port);
   NEXT_REGISTERS_reg_14_29_inst : DLH_X1 port map( G => n12012, D => N3369, Q 
                           => NEXT_REGISTERS_14_29_port);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => N1139, CK => CLK, Q => 
                           n_1482, QN => n931_port);
   NEXT_REGISTERS_reg_14_28_inst : DLH_X1 port map( G => n12012, D => N3368, Q 
                           => NEXT_REGISTERS_14_28_port);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => N1138, CK => CLK, Q => 
                           n_1483, QN => n932_port);
   NEXT_REGISTERS_reg_14_27_inst : DLH_X1 port map( G => n12012, D => N3367, Q 
                           => NEXT_REGISTERS_14_27_port);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => N1137, CK => CLK, Q => 
                           n_1484, QN => n933_port);
   NEXT_REGISTERS_reg_14_26_inst : DLH_X1 port map( G => n12012, D => N3366, Q 
                           => NEXT_REGISTERS_14_26_port);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => N1136, CK => CLK, Q => 
                           n_1485, QN => n934_port);
   NEXT_REGISTERS_reg_14_25_inst : DLH_X1 port map( G => n12012, D => N3365, Q 
                           => NEXT_REGISTERS_14_25_port);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => N1135, CK => CLK, Q => 
                           n_1486, QN => n935_port);
   NEXT_REGISTERS_reg_14_24_inst : DLH_X1 port map( G => n12012, D => N3364, Q 
                           => NEXT_REGISTERS_14_24_port);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => N1134, CK => CLK, Q => 
                           n_1487, QN => n936_port);
   NEXT_REGISTERS_reg_14_23_inst : DLH_X1 port map( G => n12012, D => N3363, Q 
                           => NEXT_REGISTERS_14_23_port);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => N1133, CK => CLK, Q => 
                           n_1488, QN => n937_port);
   NEXT_REGISTERS_reg_14_22_inst : DLH_X1 port map( G => n12012, D => N3362, Q 
                           => NEXT_REGISTERS_14_22_port);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => N1132, CK => CLK, Q => 
                           n_1489, QN => n938_port);
   NEXT_REGISTERS_reg_14_21_inst : DLH_X1 port map( G => n12012, D => N3361, Q 
                           => NEXT_REGISTERS_14_21_port);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => N1131, CK => CLK, Q => 
                           n_1490, QN => n939_port);
   NEXT_REGISTERS_reg_14_20_inst : DLH_X1 port map( G => n12012, D => N3360, Q 
                           => NEXT_REGISTERS_14_20_port);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => N1130, CK => CLK, Q => 
                           n_1491, QN => n940_port);
   NEXT_REGISTERS_reg_14_19_inst : DLH_X1 port map( G => n12013, D => N3359, Q 
                           => NEXT_REGISTERS_14_19_port);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => N1129, CK => CLK, Q => 
                           n_1492, QN => n941_port);
   NEXT_REGISTERS_reg_14_18_inst : DLH_X1 port map( G => n12013, D => N3358, Q 
                           => NEXT_REGISTERS_14_18_port);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => N1128, CK => CLK, Q => 
                           n_1493, QN => n942_port);
   NEXT_REGISTERS_reg_14_17_inst : DLH_X1 port map( G => n12013, D => N3357, Q 
                           => NEXT_REGISTERS_14_17_port);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => N1127, CK => CLK, Q => 
                           n_1494, QN => n943_port);
   NEXT_REGISTERS_reg_14_16_inst : DLH_X1 port map( G => n12013, D => N3356, Q 
                           => NEXT_REGISTERS_14_16_port);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => N1126, CK => CLK, Q => 
                           n_1495, QN => n944_port);
   NEXT_REGISTERS_reg_14_15_inst : DLH_X1 port map( G => n12013, D => N3355, Q 
                           => NEXT_REGISTERS_14_15_port);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => N1125, CK => CLK, Q => 
                           n_1496, QN => n945_port);
   NEXT_REGISTERS_reg_14_14_inst : DLH_X1 port map( G => n12013, D => N3354, Q 
                           => NEXT_REGISTERS_14_14_port);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => N1124, CK => CLK, Q => 
                           n_1497, QN => n946_port);
   NEXT_REGISTERS_reg_14_13_inst : DLH_X1 port map( G => n12013, D => N3353, Q 
                           => NEXT_REGISTERS_14_13_port);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => N1123, CK => CLK, Q => 
                           n_1498, QN => n947_port);
   NEXT_REGISTERS_reg_14_12_inst : DLH_X1 port map( G => n12013, D => N3352, Q 
                           => NEXT_REGISTERS_14_12_port);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => N1122, CK => CLK, Q => 
                           n_1499, QN => n948_port);
   NEXT_REGISTERS_reg_14_11_inst : DLH_X1 port map( G => n12013, D => N3351, Q 
                           => NEXT_REGISTERS_14_11_port);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => N1121, CK => CLK, Q => 
                           n_1500, QN => n949_port);
   NEXT_REGISTERS_reg_14_10_inst : DLH_X1 port map( G => n12013, D => N3350, Q 
                           => NEXT_REGISTERS_14_10_port);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => N1120, CK => CLK, Q => 
                           n_1501, QN => n950_port);
   NEXT_REGISTERS_reg_14_9_inst : DLH_X1 port map( G => n12013, D => N3349, Q 
                           => NEXT_REGISTERS_14_9_port);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => N1119, CK => CLK, Q => 
                           n_1502, QN => n951_port);
   NEXT_REGISTERS_reg_14_8_inst : DLH_X1 port map( G => n12014, D => N3348, Q 
                           => NEXT_REGISTERS_14_8_port);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => N1118, CK => CLK, Q => 
                           n_1503, QN => n952_port);
   NEXT_REGISTERS_reg_14_7_inst : DLH_X1 port map( G => n12014, D => N3347, Q 
                           => NEXT_REGISTERS_14_7_port);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => N1117, CK => CLK, Q => 
                           n_1504, QN => n953_port);
   NEXT_REGISTERS_reg_14_6_inst : DLH_X1 port map( G => n12014, D => N3346, Q 
                           => NEXT_REGISTERS_14_6_port);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => N1116, CK => CLK, Q => 
                           n_1505, QN => n954_port);
   NEXT_REGISTERS_reg_14_5_inst : DLH_X1 port map( G => n12014, D => N3345, Q 
                           => NEXT_REGISTERS_14_5_port);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => N1115, CK => CLK, Q => 
                           n_1506, QN => n955_port);
   NEXT_REGISTERS_reg_14_4_inst : DLH_X1 port map( G => n12014, D => N3344, Q 
                           => NEXT_REGISTERS_14_4_port);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => N1114, CK => CLK, Q => 
                           n_1507, QN => n956_port);
   NEXT_REGISTERS_reg_14_3_inst : DLH_X1 port map( G => n12014, D => N3343, Q 
                           => NEXT_REGISTERS_14_3_port);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => N1113, CK => CLK, Q => 
                           n_1508, QN => n957_port);
   NEXT_REGISTERS_reg_14_2_inst : DLH_X1 port map( G => n12014, D => N3342, Q 
                           => NEXT_REGISTERS_14_2_port);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => N1112, CK => CLK, Q => 
                           n_1509, QN => n958_port);
   NEXT_REGISTERS_reg_14_1_inst : DLH_X1 port map( G => n12014, D => N3341, Q 
                           => NEXT_REGISTERS_14_1_port);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => N1111, CK => CLK, Q => 
                           n_1510, QN => n959_port);
   NEXT_REGISTERS_reg_14_0_inst : DLH_X1 port map( G => n12014, D => N3340, Q 
                           => NEXT_REGISTERS_14_0_port);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => N1110, CK => CLK, Q => 
                           n_1511, QN => n960_port);
   NEXT_REGISTERS_reg_15_63_inst : DLH_X1 port map( G => n12018, D => N3338, Q 
                           => NEXT_REGISTERS_15_63_port);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => N1109, CK => CLK, Q => 
                           n10541, QN => n961_port);
   NEXT_REGISTERS_reg_15_62_inst : DLH_X1 port map( G => n12018, D => N3337, Q 
                           => NEXT_REGISTERS_15_62_port);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => N1108, CK => CLK, Q => 
                           n10539, QN => n962_port);
   NEXT_REGISTERS_reg_15_61_inst : DLH_X1 port map( G => n12018, D => N3336, Q 
                           => NEXT_REGISTERS_15_61_port);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => N1107, CK => CLK, Q => 
                           n10537, QN => n963_port);
   NEXT_REGISTERS_reg_15_60_inst : DLH_X1 port map( G => n12018, D => N3335, Q 
                           => NEXT_REGISTERS_15_60_port);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => N1106, CK => CLK, Q => 
                           n10535, QN => n964_port);
   NEXT_REGISTERS_reg_15_59_inst : DLH_X1 port map( G => n12018, D => N3334, Q 
                           => NEXT_REGISTERS_15_59_port);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => N1105, CK => CLK, Q => 
                           n10533, QN => n965_port);
   NEXT_REGISTERS_reg_15_58_inst : DLH_X1 port map( G => n12018, D => N3333, Q 
                           => NEXT_REGISTERS_15_58_port);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => N1104, CK => CLK, Q => 
                           n10531, QN => n966_port);
   NEXT_REGISTERS_reg_15_57_inst : DLH_X1 port map( G => n12018, D => N3332, Q 
                           => NEXT_REGISTERS_15_57_port);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => N1103, CK => CLK, Q => 
                           n10529, QN => n967_port);
   NEXT_REGISTERS_reg_15_56_inst : DLH_X1 port map( G => n12018, D => N3331, Q 
                           => NEXT_REGISTERS_15_56_port);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => N1102, CK => CLK, Q => 
                           n10527, QN => n968_port);
   NEXT_REGISTERS_reg_15_55_inst : DLH_X1 port map( G => n12018, D => N3330, Q 
                           => NEXT_REGISTERS_15_55_port);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => N1101, CK => CLK, Q => 
                           n10525, QN => n969_port);
   NEXT_REGISTERS_reg_15_54_inst : DLH_X1 port map( G => n12018, D => N3329, Q 
                           => NEXT_REGISTERS_15_54_port);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => N1100, CK => CLK, Q => 
                           n10523, QN => n970_port);
   NEXT_REGISTERS_reg_15_53_inst : DLH_X1 port map( G => n12018, D => N3328, Q 
                           => NEXT_REGISTERS_15_53_port);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => N1099, CK => CLK, Q => 
                           n10521, QN => n971_port);
   NEXT_REGISTERS_reg_15_52_inst : DLH_X1 port map( G => n12019, D => N3327, Q 
                           => NEXT_REGISTERS_15_52_port);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => N1098, CK => CLK, Q => 
                           n10519, QN => n972_port);
   NEXT_REGISTERS_reg_15_51_inst : DLH_X1 port map( G => n12019, D => N3326, Q 
                           => NEXT_REGISTERS_15_51_port);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => N1097, CK => CLK, Q => 
                           n10517, QN => n973_port);
   NEXT_REGISTERS_reg_15_50_inst : DLH_X1 port map( G => n12019, D => N3325, Q 
                           => NEXT_REGISTERS_15_50_port);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => N1096, CK => CLK, Q => 
                           n10515, QN => n974_port);
   NEXT_REGISTERS_reg_15_49_inst : DLH_X1 port map( G => n12019, D => N3324, Q 
                           => NEXT_REGISTERS_15_49_port);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => N1095, CK => CLK, Q => 
                           n10513, QN => n975_port);
   NEXT_REGISTERS_reg_15_48_inst : DLH_X1 port map( G => n12019, D => N3323, Q 
                           => NEXT_REGISTERS_15_48_port);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => N1094, CK => CLK, Q => 
                           n10511, QN => n976_port);
   NEXT_REGISTERS_reg_15_47_inst : DLH_X1 port map( G => n12019, D => N3322, Q 
                           => NEXT_REGISTERS_15_47_port);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => N1093, CK => CLK, Q => 
                           n10509, QN => n977_port);
   NEXT_REGISTERS_reg_15_46_inst : DLH_X1 port map( G => n12019, D => N3321, Q 
                           => NEXT_REGISTERS_15_46_port);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => N1092, CK => CLK, Q => 
                           n10507, QN => n978_port);
   NEXT_REGISTERS_reg_15_45_inst : DLH_X1 port map( G => n12019, D => N3320, Q 
                           => NEXT_REGISTERS_15_45_port);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => N1091, CK => CLK, Q => 
                           n10505, QN => n979_port);
   NEXT_REGISTERS_reg_15_44_inst : DLH_X1 port map( G => n12019, D => N3319, Q 
                           => NEXT_REGISTERS_15_44_port);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => N1090, CK => CLK, Q => 
                           n10503, QN => n980_port);
   NEXT_REGISTERS_reg_15_43_inst : DLH_X1 port map( G => n12019, D => N3318, Q 
                           => NEXT_REGISTERS_15_43_port);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => N1089, CK => CLK, Q => 
                           n10501, QN => n981_port);
   NEXT_REGISTERS_reg_15_42_inst : DLH_X1 port map( G => n12019, D => N3317, Q 
                           => NEXT_REGISTERS_15_42_port);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => N1088, CK => CLK, Q => 
                           n10499, QN => n982_port);
   NEXT_REGISTERS_reg_15_41_inst : DLH_X1 port map( G => n12020, D => N3316, Q 
                           => NEXT_REGISTERS_15_41_port);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => N1087, CK => CLK, Q => 
                           n10497, QN => n983_port);
   NEXT_REGISTERS_reg_15_40_inst : DLH_X1 port map( G => n12020, D => N3315, Q 
                           => NEXT_REGISTERS_15_40_port);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => N1086, CK => CLK, Q => 
                           n10495, QN => n984_port);
   NEXT_REGISTERS_reg_15_39_inst : DLH_X1 port map( G => n12020, D => N3314, Q 
                           => NEXT_REGISTERS_15_39_port);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => N1085, CK => CLK, Q => 
                           n10493, QN => n985_port);
   NEXT_REGISTERS_reg_15_38_inst : DLH_X1 port map( G => n12020, D => N3313, Q 
                           => NEXT_REGISTERS_15_38_port);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => N1084, CK => CLK, Q => 
                           n10491, QN => n986_port);
   NEXT_REGISTERS_reg_15_37_inst : DLH_X1 port map( G => n12020, D => N3312, Q 
                           => NEXT_REGISTERS_15_37_port);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => N1083, CK => CLK, Q => 
                           n10489, QN => n987_port);
   NEXT_REGISTERS_reg_15_36_inst : DLH_X1 port map( G => n12020, D => N3311, Q 
                           => NEXT_REGISTERS_15_36_port);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => N1082, CK => CLK, Q => 
                           n10487, QN => n988_port);
   NEXT_REGISTERS_reg_15_35_inst : DLH_X1 port map( G => n12020, D => N3310, Q 
                           => NEXT_REGISTERS_15_35_port);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => N1081, CK => CLK, Q => 
                           n10485, QN => n989_port);
   NEXT_REGISTERS_reg_15_34_inst : DLH_X1 port map( G => n12020, D => N3309, Q 
                           => NEXT_REGISTERS_15_34_port);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => N1080, CK => CLK, Q => 
                           n10483, QN => n990_port);
   NEXT_REGISTERS_reg_15_33_inst : DLH_X1 port map( G => n12020, D => N3308, Q 
                           => NEXT_REGISTERS_15_33_port);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => N1079, CK => CLK, Q => 
                           n10481, QN => n991_port);
   NEXT_REGISTERS_reg_15_32_inst : DLH_X1 port map( G => n12020, D => N3307, Q 
                           => NEXT_REGISTERS_15_32_port);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => N1078, CK => CLK, Q => 
                           n10479, QN => n992_port);
   NEXT_REGISTERS_reg_15_31_inst : DLH_X1 port map( G => n12020, D => N3306, Q 
                           => NEXT_REGISTERS_15_31_port);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => N1077, CK => CLK, Q => 
                           n10477, QN => n993_port);
   NEXT_REGISTERS_reg_15_30_inst : DLH_X1 port map( G => n12021, D => N3305, Q 
                           => NEXT_REGISTERS_15_30_port);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => N1076, CK => CLK, Q => 
                           n10475, QN => n994_port);
   NEXT_REGISTERS_reg_15_29_inst : DLH_X1 port map( G => n12021, D => N3304, Q 
                           => NEXT_REGISTERS_15_29_port);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => N1075, CK => CLK, Q => 
                           n10473, QN => n995_port);
   NEXT_REGISTERS_reg_15_28_inst : DLH_X1 port map( G => n12021, D => N3303, Q 
                           => NEXT_REGISTERS_15_28_port);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => N1074, CK => CLK, Q => 
                           n10471, QN => n996_port);
   NEXT_REGISTERS_reg_15_27_inst : DLH_X1 port map( G => n12021, D => N3302, Q 
                           => NEXT_REGISTERS_15_27_port);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => N1073, CK => CLK, Q => 
                           n10469, QN => n997_port);
   NEXT_REGISTERS_reg_15_26_inst : DLH_X1 port map( G => n12021, D => N3301, Q 
                           => NEXT_REGISTERS_15_26_port);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => N1072, CK => CLK, Q => 
                           n10467, QN => n998_port);
   NEXT_REGISTERS_reg_15_25_inst : DLH_X1 port map( G => n12021, D => N3300, Q 
                           => NEXT_REGISTERS_15_25_port);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => N1071, CK => CLK, Q => 
                           n10465, QN => n999_port);
   NEXT_REGISTERS_reg_15_24_inst : DLH_X1 port map( G => n12021, D => N3299, Q 
                           => NEXT_REGISTERS_15_24_port);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => N1070, CK => CLK, Q => 
                           n10463, QN => n1000_port);
   NEXT_REGISTERS_reg_15_23_inst : DLH_X1 port map( G => n12021, D => N3298, Q 
                           => NEXT_REGISTERS_15_23_port);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => N1069, CK => CLK, Q => 
                           n10461, QN => n1001_port);
   NEXT_REGISTERS_reg_15_22_inst : DLH_X1 port map( G => n12021, D => N3297, Q 
                           => NEXT_REGISTERS_15_22_port);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => N1068, CK => CLK, Q => 
                           n10459, QN => n1002_port);
   NEXT_REGISTERS_reg_15_21_inst : DLH_X1 port map( G => n12021, D => N3296, Q 
                           => NEXT_REGISTERS_15_21_port);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => N1067, CK => CLK, Q => 
                           n10457, QN => n1003_port);
   NEXT_REGISTERS_reg_15_20_inst : DLH_X1 port map( G => n12021, D => N3295, Q 
                           => NEXT_REGISTERS_15_20_port);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => N1066, CK => CLK, Q => 
                           n10455, QN => n1004_port);
   NEXT_REGISTERS_reg_15_19_inst : DLH_X1 port map( G => n12022, D => N3294, Q 
                           => NEXT_REGISTERS_15_19_port);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => N1065, CK => CLK, Q => 
                           n10453, QN => n1005_port);
   NEXT_REGISTERS_reg_15_18_inst : DLH_X1 port map( G => n12022, D => N3293, Q 
                           => NEXT_REGISTERS_15_18_port);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => N1064, CK => CLK, Q => 
                           n10451, QN => n1006_port);
   NEXT_REGISTERS_reg_15_17_inst : DLH_X1 port map( G => n12022, D => N3292, Q 
                           => NEXT_REGISTERS_15_17_port);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => N1063, CK => CLK, Q => 
                           n10449, QN => n1007_port);
   NEXT_REGISTERS_reg_15_16_inst : DLH_X1 port map( G => n12022, D => N3291, Q 
                           => NEXT_REGISTERS_15_16_port);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => N1062, CK => CLK, Q => 
                           n10447, QN => n1008_port);
   NEXT_REGISTERS_reg_15_15_inst : DLH_X1 port map( G => n12022, D => N3290, Q 
                           => NEXT_REGISTERS_15_15_port);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => N1061, CK => CLK, Q => 
                           n10445, QN => n1009_port);
   NEXT_REGISTERS_reg_15_14_inst : DLH_X1 port map( G => n12022, D => N3289, Q 
                           => NEXT_REGISTERS_15_14_port);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => N1060, CK => CLK, Q => 
                           n10443, QN => n1010_port);
   NEXT_REGISTERS_reg_15_13_inst : DLH_X1 port map( G => n12022, D => N3288, Q 
                           => NEXT_REGISTERS_15_13_port);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => N1059, CK => CLK, Q => 
                           n10441, QN => n1011_port);
   NEXT_REGISTERS_reg_15_12_inst : DLH_X1 port map( G => n12022, D => N3287, Q 
                           => NEXT_REGISTERS_15_12_port);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => N1058, CK => CLK, Q => 
                           n10439, QN => n1012_port);
   NEXT_REGISTERS_reg_15_11_inst : DLH_X1 port map( G => n12022, D => N3286, Q 
                           => NEXT_REGISTERS_15_11_port);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => N1057, CK => CLK, Q => 
                           n10437, QN => n1013_port);
   NEXT_REGISTERS_reg_15_10_inst : DLH_X1 port map( G => n12022, D => N3285, Q 
                           => NEXT_REGISTERS_15_10_port);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => N1056, CK => CLK, Q => 
                           n10435, QN => n1014_port);
   NEXT_REGISTERS_reg_15_9_inst : DLH_X1 port map( G => n12022, D => N3284, Q 
                           => NEXT_REGISTERS_15_9_port);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => N1055, CK => CLK, Q => 
                           n10433, QN => n1015_port);
   NEXT_REGISTERS_reg_15_8_inst : DLH_X1 port map( G => n12023, D => N3283, Q 
                           => NEXT_REGISTERS_15_8_port);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => N1054, CK => CLK, Q => 
                           n10431, QN => n1016_port);
   NEXT_REGISTERS_reg_15_7_inst : DLH_X1 port map( G => n12023, D => N3282, Q 
                           => NEXT_REGISTERS_15_7_port);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => N1053, CK => CLK, Q => 
                           n10429, QN => n1017_port);
   NEXT_REGISTERS_reg_15_6_inst : DLH_X1 port map( G => n12023, D => N3281, Q 
                           => NEXT_REGISTERS_15_6_port);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => N1052, CK => CLK, Q => 
                           n10427, QN => n1018_port);
   NEXT_REGISTERS_reg_15_5_inst : DLH_X1 port map( G => n12023, D => N3280, Q 
                           => NEXT_REGISTERS_15_5_port);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => N1051, CK => CLK, Q => 
                           n10425, QN => n1019_port);
   NEXT_REGISTERS_reg_15_4_inst : DLH_X1 port map( G => n12023, D => N3279, Q 
                           => NEXT_REGISTERS_15_4_port);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => N1050, CK => CLK, Q => 
                           n10423, QN => n1020_port);
   NEXT_REGISTERS_reg_15_3_inst : DLH_X1 port map( G => n12023, D => N3278, Q 
                           => NEXT_REGISTERS_15_3_port);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => N1049, CK => CLK, Q => 
                           n10421, QN => n1021_port);
   NEXT_REGISTERS_reg_15_2_inst : DLH_X1 port map( G => n12023, D => N3277, Q 
                           => NEXT_REGISTERS_15_2_port);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => N1048, CK => CLK, Q => 
                           n10419, QN => n1022_port);
   NEXT_REGISTERS_reg_15_1_inst : DLH_X1 port map( G => n12023, D => N3276, Q 
                           => NEXT_REGISTERS_15_1_port);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => N1047, CK => CLK, Q => 
                           n10417, QN => n1023_port);
   NEXT_REGISTERS_reg_15_0_inst : DLH_X1 port map( G => n12023, D => N3275, Q 
                           => NEXT_REGISTERS_15_0_port);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => N1046, CK => CLK, Q => 
                           n10415, QN => n1024_port);
   NEXT_REGISTERS_reg_16_63_inst : DLH_X1 port map( G => n12027, D => N3273, Q 
                           => NEXT_REGISTERS_16_63_port);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => N1045, CK => CLK, Q => 
                           n_1512, QN => n1025_port);
   NEXT_REGISTERS_reg_16_62_inst : DLH_X1 port map( G => n12027, D => N3272, Q 
                           => NEXT_REGISTERS_16_62_port);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => N1044, CK => CLK, Q => 
                           n_1513, QN => n1026_port);
   NEXT_REGISTERS_reg_16_61_inst : DLH_X1 port map( G => n12027, D => N3271, Q 
                           => NEXT_REGISTERS_16_61_port);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => N1043, CK => CLK, Q => 
                           n_1514, QN => n1027_port);
   NEXT_REGISTERS_reg_16_60_inst : DLH_X1 port map( G => n12027, D => N3270, Q 
                           => NEXT_REGISTERS_16_60_port);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => N1042, CK => CLK, Q => 
                           n_1515, QN => n1028_port);
   NEXT_REGISTERS_reg_16_59_inst : DLH_X1 port map( G => n12027, D => N3269, Q 
                           => NEXT_REGISTERS_16_59_port);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => N1041, CK => CLK, Q => 
                           n_1516, QN => n1029_port);
   NEXT_REGISTERS_reg_16_58_inst : DLH_X1 port map( G => n12027, D => N3268, Q 
                           => NEXT_REGISTERS_16_58_port);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => N1040, CK => CLK, Q => 
                           n_1517, QN => n1030_port);
   NEXT_REGISTERS_reg_16_57_inst : DLH_X1 port map( G => n12027, D => N3267, Q 
                           => NEXT_REGISTERS_16_57_port);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => N1039, CK => CLK, Q => 
                           n_1518, QN => n1031_port);
   NEXT_REGISTERS_reg_16_56_inst : DLH_X1 port map( G => n12027, D => N3266, Q 
                           => NEXT_REGISTERS_16_56_port);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => N1038, CK => CLK, Q => 
                           n_1519, QN => n1032_port);
   NEXT_REGISTERS_reg_16_55_inst : DLH_X1 port map( G => n12027, D => N3265, Q 
                           => NEXT_REGISTERS_16_55_port);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => N1037, CK => CLK, Q => 
                           n_1520, QN => n1033_port);
   NEXT_REGISTERS_reg_16_54_inst : DLH_X1 port map( G => n12027, D => N3264, Q 
                           => NEXT_REGISTERS_16_54_port);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => N1036, CK => CLK, Q => 
                           n_1521, QN => n1034_port);
   NEXT_REGISTERS_reg_16_53_inst : DLH_X1 port map( G => n12027, D => N3263, Q 
                           => NEXT_REGISTERS_16_53_port);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => N1035, CK => CLK, Q => 
                           n_1522, QN => n1035_port);
   NEXT_REGISTERS_reg_16_52_inst : DLH_X1 port map( G => n12028, D => N3262, Q 
                           => NEXT_REGISTERS_16_52_port);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => N1034, CK => CLK, Q => 
                           n_1523, QN => n1036_port);
   NEXT_REGISTERS_reg_16_51_inst : DLH_X1 port map( G => n12028, D => N3261, Q 
                           => NEXT_REGISTERS_16_51_port);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => N1033, CK => CLK, Q => 
                           n_1524, QN => n1037_port);
   NEXT_REGISTERS_reg_16_50_inst : DLH_X1 port map( G => n12028, D => N3260, Q 
                           => NEXT_REGISTERS_16_50_port);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => N1032, CK => CLK, Q => 
                           n_1525, QN => n1038_port);
   NEXT_REGISTERS_reg_16_49_inst : DLH_X1 port map( G => n12028, D => N3259, Q 
                           => NEXT_REGISTERS_16_49_port);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => N1031, CK => CLK, Q => 
                           n_1526, QN => n1039_port);
   NEXT_REGISTERS_reg_16_48_inst : DLH_X1 port map( G => n12028, D => N3258, Q 
                           => NEXT_REGISTERS_16_48_port);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => N1030, CK => CLK, Q => 
                           n_1527, QN => n1040_port);
   NEXT_REGISTERS_reg_16_47_inst : DLH_X1 port map( G => n12028, D => N3257, Q 
                           => NEXT_REGISTERS_16_47_port);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => N1029, CK => CLK, Q => 
                           n_1528, QN => n1041_port);
   NEXT_REGISTERS_reg_16_46_inst : DLH_X1 port map( G => n12028, D => N3256, Q 
                           => NEXT_REGISTERS_16_46_port);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => N1028, CK => CLK, Q => 
                           n_1529, QN => n1042_port);
   NEXT_REGISTERS_reg_16_45_inst : DLH_X1 port map( G => n12028, D => N3255, Q 
                           => NEXT_REGISTERS_16_45_port);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => N1027, CK => CLK, Q => 
                           n_1530, QN => n1043_port);
   NEXT_REGISTERS_reg_16_44_inst : DLH_X1 port map( G => n12028, D => N3254, Q 
                           => NEXT_REGISTERS_16_44_port);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => N1026, CK => CLK, Q => 
                           n_1531, QN => n1044_port);
   NEXT_REGISTERS_reg_16_43_inst : DLH_X1 port map( G => n12028, D => N3253, Q 
                           => NEXT_REGISTERS_16_43_port);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => N1025, CK => CLK, Q => 
                           n_1532, QN => n1045_port);
   NEXT_REGISTERS_reg_16_42_inst : DLH_X1 port map( G => n12028, D => N3252, Q 
                           => NEXT_REGISTERS_16_42_port);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => N1024, CK => CLK, Q => 
                           n_1533, QN => n1046_port);
   NEXT_REGISTERS_reg_16_41_inst : DLH_X1 port map( G => n12029, D => N3251, Q 
                           => NEXT_REGISTERS_16_41_port);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => N1023, CK => CLK, Q => 
                           n_1534, QN => n1047_port);
   NEXT_REGISTERS_reg_16_40_inst : DLH_X1 port map( G => n12029, D => N3250, Q 
                           => NEXT_REGISTERS_16_40_port);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => N1022, CK => CLK, Q => 
                           n_1535, QN => n1048_port);
   NEXT_REGISTERS_reg_16_39_inst : DLH_X1 port map( G => n12029, D => N3249, Q 
                           => NEXT_REGISTERS_16_39_port);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => N1021, CK => CLK, Q => 
                           n_1536, QN => n1049_port);
   NEXT_REGISTERS_reg_16_38_inst : DLH_X1 port map( G => n12029, D => N3248, Q 
                           => NEXT_REGISTERS_16_38_port);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => N1020, CK => CLK, Q => 
                           n_1537, QN => n1050_port);
   NEXT_REGISTERS_reg_16_37_inst : DLH_X1 port map( G => n12029, D => N3247, Q 
                           => NEXT_REGISTERS_16_37_port);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => N1019, CK => CLK, Q => 
                           n_1538, QN => n1051_port);
   NEXT_REGISTERS_reg_16_36_inst : DLH_X1 port map( G => n12029, D => N3246, Q 
                           => NEXT_REGISTERS_16_36_port);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => N1018, CK => CLK, Q => 
                           n_1539, QN => n1052_port);
   NEXT_REGISTERS_reg_16_35_inst : DLH_X1 port map( G => n12029, D => N3245, Q 
                           => NEXT_REGISTERS_16_35_port);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => N1017, CK => CLK, Q => 
                           n_1540, QN => n1053_port);
   NEXT_REGISTERS_reg_16_34_inst : DLH_X1 port map( G => n12029, D => N3244, Q 
                           => NEXT_REGISTERS_16_34_port);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => N1016, CK => CLK, Q => 
                           n_1541, QN => n1054_port);
   NEXT_REGISTERS_reg_16_33_inst : DLH_X1 port map( G => n12029, D => N3243, Q 
                           => NEXT_REGISTERS_16_33_port);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => N1015, CK => CLK, Q => 
                           n_1542, QN => n1055_port);
   NEXT_REGISTERS_reg_16_32_inst : DLH_X1 port map( G => n12029, D => N3242, Q 
                           => NEXT_REGISTERS_16_32_port);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => N1014, CK => CLK, Q => 
                           n_1543, QN => n1056_port);
   NEXT_REGISTERS_reg_16_31_inst : DLH_X1 port map( G => n12029, D => N3241, Q 
                           => NEXT_REGISTERS_16_31_port);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => N1013, CK => CLK, Q => 
                           n_1544, QN => n1057_port);
   NEXT_REGISTERS_reg_16_30_inst : DLH_X1 port map( G => n12030, D => N3240, Q 
                           => NEXT_REGISTERS_16_30_port);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => N1012, CK => CLK, Q => 
                           n_1545, QN => n1058_port);
   NEXT_REGISTERS_reg_16_29_inst : DLH_X1 port map( G => n12030, D => N3239, Q 
                           => NEXT_REGISTERS_16_29_port);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => N1011, CK => CLK, Q => 
                           n_1546, QN => n1059_port);
   NEXT_REGISTERS_reg_16_28_inst : DLH_X1 port map( G => n12030, D => N3238, Q 
                           => NEXT_REGISTERS_16_28_port);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => N1010, CK => CLK, Q => 
                           n_1547, QN => n1060_port);
   NEXT_REGISTERS_reg_16_27_inst : DLH_X1 port map( G => n12030, D => N3237, Q 
                           => NEXT_REGISTERS_16_27_port);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => N1009, CK => CLK, Q => 
                           n_1548, QN => n1061_port);
   NEXT_REGISTERS_reg_16_26_inst : DLH_X1 port map( G => n12030, D => N3236, Q 
                           => NEXT_REGISTERS_16_26_port);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => N1008, CK => CLK, Q => 
                           n_1549, QN => n1062_port);
   NEXT_REGISTERS_reg_16_25_inst : DLH_X1 port map( G => n12030, D => N3235, Q 
                           => NEXT_REGISTERS_16_25_port);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => N1007, CK => CLK, Q => 
                           n_1550, QN => n1063_port);
   NEXT_REGISTERS_reg_16_24_inst : DLH_X1 port map( G => n12030, D => N3234, Q 
                           => NEXT_REGISTERS_16_24_port);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => N1006, CK => CLK, Q => 
                           n_1551, QN => n1064_port);
   NEXT_REGISTERS_reg_16_23_inst : DLH_X1 port map( G => n12030, D => N3233, Q 
                           => NEXT_REGISTERS_16_23_port);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => N1005, CK => CLK, Q => 
                           n_1552, QN => n1065_port);
   NEXT_REGISTERS_reg_16_22_inst : DLH_X1 port map( G => n12030, D => N3232, Q 
                           => NEXT_REGISTERS_16_22_port);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => N1004, CK => CLK, Q => 
                           n_1553, QN => n1066_port);
   NEXT_REGISTERS_reg_16_21_inst : DLH_X1 port map( G => n12030, D => N3231, Q 
                           => NEXT_REGISTERS_16_21_port);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => N1003, CK => CLK, Q => 
                           n_1554, QN => n1067_port);
   NEXT_REGISTERS_reg_16_20_inst : DLH_X1 port map( G => n12030, D => N3230, Q 
                           => NEXT_REGISTERS_16_20_port);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => N1002, CK => CLK, Q => 
                           n_1555, QN => n1068_port);
   NEXT_REGISTERS_reg_16_19_inst : DLH_X1 port map( G => n12031, D => N3229, Q 
                           => NEXT_REGISTERS_16_19_port);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => N1001, CK => CLK, Q => 
                           n_1556, QN => n1069_port);
   NEXT_REGISTERS_reg_16_18_inst : DLH_X1 port map( G => n12031, D => N3228, Q 
                           => NEXT_REGISTERS_16_18_port);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => N1000, CK => CLK, Q => 
                           n_1557, QN => n1070_port);
   NEXT_REGISTERS_reg_16_17_inst : DLH_X1 port map( G => n12031, D => N3227, Q 
                           => NEXT_REGISTERS_16_17_port);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => N999, CK => CLK, Q => 
                           n_1558, QN => n1071_port);
   NEXT_REGISTERS_reg_16_16_inst : DLH_X1 port map( G => n12031, D => N3226, Q 
                           => NEXT_REGISTERS_16_16_port);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => N998, CK => CLK, Q => 
                           n_1559, QN => n1072_port);
   NEXT_REGISTERS_reg_16_15_inst : DLH_X1 port map( G => n12031, D => N3225, Q 
                           => NEXT_REGISTERS_16_15_port);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => N997, CK => CLK, Q => 
                           n_1560, QN => n1073_port);
   NEXT_REGISTERS_reg_16_14_inst : DLH_X1 port map( G => n12031, D => N3224, Q 
                           => NEXT_REGISTERS_16_14_port);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => N996, CK => CLK, Q => 
                           n_1561, QN => n1074_port);
   NEXT_REGISTERS_reg_16_13_inst : DLH_X1 port map( G => n12031, D => N3223, Q 
                           => NEXT_REGISTERS_16_13_port);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => N995, CK => CLK, Q => 
                           n_1562, QN => n1075_port);
   NEXT_REGISTERS_reg_16_12_inst : DLH_X1 port map( G => n12031, D => N3222, Q 
                           => NEXT_REGISTERS_16_12_port);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => N994, CK => CLK, Q => 
                           n_1563, QN => n1076_port);
   NEXT_REGISTERS_reg_16_11_inst : DLH_X1 port map( G => n12031, D => N3221, Q 
                           => NEXT_REGISTERS_16_11_port);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => N993, CK => CLK, Q => 
                           n_1564, QN => n1077_port);
   NEXT_REGISTERS_reg_16_10_inst : DLH_X1 port map( G => n12031, D => N3220, Q 
                           => NEXT_REGISTERS_16_10_port);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => N992, CK => CLK, Q => 
                           n_1565, QN => n1078_port);
   NEXT_REGISTERS_reg_16_9_inst : DLH_X1 port map( G => n12031, D => N3219, Q 
                           => NEXT_REGISTERS_16_9_port);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => N991, CK => CLK, Q => n_1566
                           , QN => n1079_port);
   NEXT_REGISTERS_reg_16_8_inst : DLH_X1 port map( G => n12032, D => N3218, Q 
                           => NEXT_REGISTERS_16_8_port);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => N990, CK => CLK, Q => n_1567
                           , QN => n1080_port);
   NEXT_REGISTERS_reg_16_7_inst : DLH_X1 port map( G => n12032, D => N3217, Q 
                           => NEXT_REGISTERS_16_7_port);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => N989, CK => CLK, Q => n_1568
                           , QN => n1081_port);
   NEXT_REGISTERS_reg_16_6_inst : DLH_X1 port map( G => n12032, D => N3216, Q 
                           => NEXT_REGISTERS_16_6_port);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => N988, CK => CLK, Q => n_1569
                           , QN => n1082_port);
   NEXT_REGISTERS_reg_16_5_inst : DLH_X1 port map( G => n12032, D => N3215, Q 
                           => NEXT_REGISTERS_16_5_port);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => N987, CK => CLK, Q => n_1570
                           , QN => n1083_port);
   NEXT_REGISTERS_reg_16_4_inst : DLH_X1 port map( G => n12032, D => N3214, Q 
                           => NEXT_REGISTERS_16_4_port);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => N986, CK => CLK, Q => n_1571
                           , QN => n1084_port);
   NEXT_REGISTERS_reg_16_3_inst : DLH_X1 port map( G => n12032, D => N3213, Q 
                           => NEXT_REGISTERS_16_3_port);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => N985, CK => CLK, Q => n_1572
                           , QN => n1085_port);
   NEXT_REGISTERS_reg_16_2_inst : DLH_X1 port map( G => n12032, D => N3212, Q 
                           => NEXT_REGISTERS_16_2_port);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => N984, CK => CLK, Q => n_1573
                           , QN => n1086_port);
   NEXT_REGISTERS_reg_16_1_inst : DLH_X1 port map( G => n12032, D => N3211, Q 
                           => NEXT_REGISTERS_16_1_port);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => N983, CK => CLK, Q => n_1574
                           , QN => n1087_port);
   NEXT_REGISTERS_reg_16_0_inst : DLH_X1 port map( G => n12032, D => N3210, Q 
                           => NEXT_REGISTERS_16_0_port);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => N982, CK => CLK, Q => n_1575
                           , QN => n1088_port);
   NEXT_REGISTERS_reg_17_63_inst : DLH_X1 port map( G => n12036, D => N3208, Q 
                           => NEXT_REGISTERS_17_63_port);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => N981, CK => CLK, Q => 
                           n_1576, QN => n1089_port);
   NEXT_REGISTERS_reg_17_62_inst : DLH_X1 port map( G => n12036, D => N3207, Q 
                           => NEXT_REGISTERS_17_62_port);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => N980, CK => CLK, Q => 
                           n_1577, QN => n1090_port);
   NEXT_REGISTERS_reg_17_61_inst : DLH_X1 port map( G => n12036, D => N3206, Q 
                           => NEXT_REGISTERS_17_61_port);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => N979, CK => CLK, Q => 
                           n_1578, QN => n1091_port);
   NEXT_REGISTERS_reg_17_60_inst : DLH_X1 port map( G => n12036, D => N3205, Q 
                           => NEXT_REGISTERS_17_60_port);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => N978, CK => CLK, Q => 
                           n_1579, QN => n1092_port);
   NEXT_REGISTERS_reg_17_59_inst : DLH_X1 port map( G => n12036, D => N3204, Q 
                           => NEXT_REGISTERS_17_59_port);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => N977, CK => CLK, Q => 
                           n_1580, QN => n1093_port);
   NEXT_REGISTERS_reg_17_58_inst : DLH_X1 port map( G => n12036, D => N3203, Q 
                           => NEXT_REGISTERS_17_58_port);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => N976, CK => CLK, Q => 
                           n_1581, QN => n1094_port);
   NEXT_REGISTERS_reg_17_57_inst : DLH_X1 port map( G => n12036, D => N3202, Q 
                           => NEXT_REGISTERS_17_57_port);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => N975, CK => CLK, Q => 
                           n_1582, QN => n1095_port);
   NEXT_REGISTERS_reg_17_56_inst : DLH_X1 port map( G => n12036, D => N3201, Q 
                           => NEXT_REGISTERS_17_56_port);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => N974, CK => CLK, Q => 
                           n_1583, QN => n1096_port);
   NEXT_REGISTERS_reg_17_55_inst : DLH_X1 port map( G => n12036, D => N3200, Q 
                           => NEXT_REGISTERS_17_55_port);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => N973, CK => CLK, Q => 
                           n_1584, QN => n1097_port);
   NEXT_REGISTERS_reg_17_54_inst : DLH_X1 port map( G => n12036, D => N3199, Q 
                           => NEXT_REGISTERS_17_54_port);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => N972, CK => CLK, Q => 
                           n_1585, QN => n1098_port);
   NEXT_REGISTERS_reg_17_53_inst : DLH_X1 port map( G => n12036, D => N3198, Q 
                           => NEXT_REGISTERS_17_53_port);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => N971, CK => CLK, Q => 
                           n_1586, QN => n1099_port);
   NEXT_REGISTERS_reg_17_52_inst : DLH_X1 port map( G => n12037, D => N3197, Q 
                           => NEXT_REGISTERS_17_52_port);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => N970, CK => CLK, Q => 
                           n_1587, QN => n1100_port);
   NEXT_REGISTERS_reg_17_51_inst : DLH_X1 port map( G => n12037, D => N3196, Q 
                           => NEXT_REGISTERS_17_51_port);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => N969, CK => CLK, Q => 
                           n_1588, QN => n1101_port);
   NEXT_REGISTERS_reg_17_50_inst : DLH_X1 port map( G => n12037, D => N3195, Q 
                           => NEXT_REGISTERS_17_50_port);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => N968, CK => CLK, Q => 
                           n_1589, QN => n1102_port);
   NEXT_REGISTERS_reg_17_49_inst : DLH_X1 port map( G => n12037, D => N3194, Q 
                           => NEXT_REGISTERS_17_49_port);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => N967, CK => CLK, Q => 
                           n_1590, QN => n1103_port);
   NEXT_REGISTERS_reg_17_48_inst : DLH_X1 port map( G => n12037, D => N3193, Q 
                           => NEXT_REGISTERS_17_48_port);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => N966, CK => CLK, Q => 
                           n_1591, QN => n1104_port);
   NEXT_REGISTERS_reg_17_47_inst : DLH_X1 port map( G => n12037, D => N3192, Q 
                           => NEXT_REGISTERS_17_47_port);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => N965, CK => CLK, Q => 
                           n_1592, QN => n1105_port);
   NEXT_REGISTERS_reg_17_46_inst : DLH_X1 port map( G => n12037, D => N3191, Q 
                           => NEXT_REGISTERS_17_46_port);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => N964, CK => CLK, Q => 
                           n_1593, QN => n1106_port);
   NEXT_REGISTERS_reg_17_45_inst : DLH_X1 port map( G => n12037, D => N3190, Q 
                           => NEXT_REGISTERS_17_45_port);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => N963, CK => CLK, Q => 
                           n_1594, QN => n1107_port);
   NEXT_REGISTERS_reg_17_44_inst : DLH_X1 port map( G => n12037, D => N3189, Q 
                           => NEXT_REGISTERS_17_44_port);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => N962, CK => CLK, Q => 
                           n_1595, QN => n1108_port);
   NEXT_REGISTERS_reg_17_43_inst : DLH_X1 port map( G => n12037, D => N3188, Q 
                           => NEXT_REGISTERS_17_43_port);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => N961, CK => CLK, Q => 
                           n_1596, QN => n1109_port);
   NEXT_REGISTERS_reg_17_42_inst : DLH_X1 port map( G => n12037, D => N3187, Q 
                           => NEXT_REGISTERS_17_42_port);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => N960, CK => CLK, Q => 
                           n_1597, QN => n1110_port);
   NEXT_REGISTERS_reg_17_41_inst : DLH_X1 port map( G => n12038, D => N3186, Q 
                           => NEXT_REGISTERS_17_41_port);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => N959, CK => CLK, Q => 
                           n_1598, QN => n1111_port);
   NEXT_REGISTERS_reg_17_40_inst : DLH_X1 port map( G => n12038, D => N3185, Q 
                           => NEXT_REGISTERS_17_40_port);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => N958, CK => CLK, Q => 
                           n_1599, QN => n1112_port);
   NEXT_REGISTERS_reg_17_39_inst : DLH_X1 port map( G => n12038, D => N3184, Q 
                           => NEXT_REGISTERS_17_39_port);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => N957, CK => CLK, Q => 
                           n_1600, QN => n1113_port);
   NEXT_REGISTERS_reg_17_38_inst : DLH_X1 port map( G => n12038, D => N3183, Q 
                           => NEXT_REGISTERS_17_38_port);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => N956, CK => CLK, Q => 
                           n_1601, QN => n1114_port);
   NEXT_REGISTERS_reg_17_37_inst : DLH_X1 port map( G => n12038, D => N3182, Q 
                           => NEXT_REGISTERS_17_37_port);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => N955, CK => CLK, Q => 
                           n_1602, QN => n1115_port);
   NEXT_REGISTERS_reg_17_36_inst : DLH_X1 port map( G => n12038, D => N3181, Q 
                           => NEXT_REGISTERS_17_36_port);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => N954, CK => CLK, Q => 
                           n_1603, QN => n1116_port);
   NEXT_REGISTERS_reg_17_35_inst : DLH_X1 port map( G => n12038, D => N3180, Q 
                           => NEXT_REGISTERS_17_35_port);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => N953, CK => CLK, Q => 
                           n_1604, QN => n1117_port);
   NEXT_REGISTERS_reg_17_34_inst : DLH_X1 port map( G => n12038, D => N3179, Q 
                           => NEXT_REGISTERS_17_34_port);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => N952, CK => CLK, Q => 
                           n_1605, QN => n1118_port);
   NEXT_REGISTERS_reg_17_33_inst : DLH_X1 port map( G => n12038, D => N3178, Q 
                           => NEXT_REGISTERS_17_33_port);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => N951, CK => CLK, Q => 
                           n_1606, QN => n1119_port);
   NEXT_REGISTERS_reg_17_32_inst : DLH_X1 port map( G => n12038, D => N3177, Q 
                           => NEXT_REGISTERS_17_32_port);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => N950, CK => CLK, Q => 
                           n_1607, QN => n1120_port);
   NEXT_REGISTERS_reg_17_31_inst : DLH_X1 port map( G => n12038, D => N3176, Q 
                           => NEXT_REGISTERS_17_31_port);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => N949, CK => CLK, Q => 
                           n_1608, QN => n1121_port);
   NEXT_REGISTERS_reg_17_30_inst : DLH_X1 port map( G => n12039, D => N3175, Q 
                           => NEXT_REGISTERS_17_30_port);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => N948, CK => CLK, Q => 
                           n_1609, QN => n1122_port);
   NEXT_REGISTERS_reg_17_29_inst : DLH_X1 port map( G => n12039, D => N3174, Q 
                           => NEXT_REGISTERS_17_29_port);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => N947, CK => CLK, Q => 
                           n_1610, QN => n1123_port);
   NEXT_REGISTERS_reg_17_28_inst : DLH_X1 port map( G => n12039, D => N3173, Q 
                           => NEXT_REGISTERS_17_28_port);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => N946, CK => CLK, Q => 
                           n_1611, QN => n1124_port);
   NEXT_REGISTERS_reg_17_27_inst : DLH_X1 port map( G => n12039, D => N3172, Q 
                           => NEXT_REGISTERS_17_27_port);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => N945, CK => CLK, Q => 
                           n_1612, QN => n1125_port);
   NEXT_REGISTERS_reg_17_26_inst : DLH_X1 port map( G => n12039, D => N3171, Q 
                           => NEXT_REGISTERS_17_26_port);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => N944, CK => CLK, Q => 
                           n_1613, QN => n1126_port);
   NEXT_REGISTERS_reg_17_25_inst : DLH_X1 port map( G => n12039, D => N3170, Q 
                           => NEXT_REGISTERS_17_25_port);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => N943, CK => CLK, Q => 
                           n_1614, QN => n1127_port);
   NEXT_REGISTERS_reg_17_24_inst : DLH_X1 port map( G => n12039, D => N3169, Q 
                           => NEXT_REGISTERS_17_24_port);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => N942, CK => CLK, Q => 
                           n_1615, QN => n1128_port);
   NEXT_REGISTERS_reg_17_23_inst : DLH_X1 port map( G => n12039, D => N3168, Q 
                           => NEXT_REGISTERS_17_23_port);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => N941, CK => CLK, Q => 
                           n_1616, QN => n1129_port);
   NEXT_REGISTERS_reg_17_22_inst : DLH_X1 port map( G => n12039, D => N3167, Q 
                           => NEXT_REGISTERS_17_22_port);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => N940, CK => CLK, Q => 
                           n_1617, QN => n1130_port);
   NEXT_REGISTERS_reg_17_21_inst : DLH_X1 port map( G => n12039, D => N3166, Q 
                           => NEXT_REGISTERS_17_21_port);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => N939, CK => CLK, Q => 
                           n_1618, QN => n1131_port);
   NEXT_REGISTERS_reg_17_20_inst : DLH_X1 port map( G => n12039, D => N3165, Q 
                           => NEXT_REGISTERS_17_20_port);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => N938, CK => CLK, Q => 
                           n_1619, QN => n1132_port);
   NEXT_REGISTERS_reg_17_19_inst : DLH_X1 port map( G => n12040, D => N3164, Q 
                           => NEXT_REGISTERS_17_19_port);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => N937, CK => CLK, Q => 
                           n_1620, QN => n1133_port);
   NEXT_REGISTERS_reg_17_18_inst : DLH_X1 port map( G => n12040, D => N3163, Q 
                           => NEXT_REGISTERS_17_18_port);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => N936, CK => CLK, Q => 
                           n_1621, QN => n1134_port);
   NEXT_REGISTERS_reg_17_17_inst : DLH_X1 port map( G => n12040, D => N3162, Q 
                           => NEXT_REGISTERS_17_17_port);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => N935, CK => CLK, Q => 
                           n_1622, QN => n1135_port);
   NEXT_REGISTERS_reg_17_16_inst : DLH_X1 port map( G => n12040, D => N3161, Q 
                           => NEXT_REGISTERS_17_16_port);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => N934, CK => CLK, Q => 
                           n_1623, QN => n1136_port);
   NEXT_REGISTERS_reg_17_15_inst : DLH_X1 port map( G => n12040, D => N3160, Q 
                           => NEXT_REGISTERS_17_15_port);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => N933, CK => CLK, Q => 
                           n_1624, QN => n1137_port);
   NEXT_REGISTERS_reg_17_14_inst : DLH_X1 port map( G => n12040, D => N3159, Q 
                           => NEXT_REGISTERS_17_14_port);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => N932, CK => CLK, Q => 
                           n_1625, QN => n1138_port);
   NEXT_REGISTERS_reg_17_13_inst : DLH_X1 port map( G => n12040, D => N3158, Q 
                           => NEXT_REGISTERS_17_13_port);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => N931, CK => CLK, Q => 
                           n_1626, QN => n1139_port);
   NEXT_REGISTERS_reg_17_12_inst : DLH_X1 port map( G => n12040, D => N3157, Q 
                           => NEXT_REGISTERS_17_12_port);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => N930, CK => CLK, Q => 
                           n_1627, QN => n1140_port);
   NEXT_REGISTERS_reg_17_11_inst : DLH_X1 port map( G => n12040, D => N3156, Q 
                           => NEXT_REGISTERS_17_11_port);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => N929, CK => CLK, Q => 
                           n_1628, QN => n1141_port);
   NEXT_REGISTERS_reg_17_10_inst : DLH_X1 port map( G => n12040, D => N3155, Q 
                           => NEXT_REGISTERS_17_10_port);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => N928, CK => CLK, Q => 
                           n_1629, QN => n1142_port);
   NEXT_REGISTERS_reg_17_9_inst : DLH_X1 port map( G => n12040, D => N3154, Q 
                           => NEXT_REGISTERS_17_9_port);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => N927, CK => CLK, Q => n_1630
                           , QN => n1143_port);
   NEXT_REGISTERS_reg_17_8_inst : DLH_X1 port map( G => n12041, D => N3153, Q 
                           => NEXT_REGISTERS_17_8_port);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => N926, CK => CLK, Q => n_1631
                           , QN => n1144_port);
   NEXT_REGISTERS_reg_17_7_inst : DLH_X1 port map( G => n12041, D => N3152, Q 
                           => NEXT_REGISTERS_17_7_port);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => N925, CK => CLK, Q => n_1632
                           , QN => n1145_port);
   NEXT_REGISTERS_reg_17_6_inst : DLH_X1 port map( G => n12041, D => N3151, Q 
                           => NEXT_REGISTERS_17_6_port);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => N924, CK => CLK, Q => n_1633
                           , QN => n1146_port);
   NEXT_REGISTERS_reg_17_5_inst : DLH_X1 port map( G => n12041, D => N3150, Q 
                           => NEXT_REGISTERS_17_5_port);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => N923, CK => CLK, Q => n_1634
                           , QN => n1147_port);
   NEXT_REGISTERS_reg_17_4_inst : DLH_X1 port map( G => n12041, D => N3149, Q 
                           => NEXT_REGISTERS_17_4_port);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => N922, CK => CLK, Q => n_1635
                           , QN => n1148_port);
   NEXT_REGISTERS_reg_17_3_inst : DLH_X1 port map( G => n12041, D => N3148, Q 
                           => NEXT_REGISTERS_17_3_port);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => N921, CK => CLK, Q => n_1636
                           , QN => n1149_port);
   NEXT_REGISTERS_reg_17_2_inst : DLH_X1 port map( G => n12041, D => N3147, Q 
                           => NEXT_REGISTERS_17_2_port);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => N920, CK => CLK, Q => n_1637
                           , QN => n1150_port);
   NEXT_REGISTERS_reg_17_1_inst : DLH_X1 port map( G => n12041, D => N3146, Q 
                           => NEXT_REGISTERS_17_1_port);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => N919, CK => CLK, Q => n_1638
                           , QN => n1151_port);
   NEXT_REGISTERS_reg_17_0_inst : DLH_X1 port map( G => n12041, D => N3145, Q 
                           => NEXT_REGISTERS_17_0_port);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => N918, CK => CLK, Q => n_1639
                           , QN => n1152_port);
   NEXT_REGISTERS_reg_18_63_inst : DLH_X1 port map( G => n12045, D => N3143, Q 
                           => NEXT_REGISTERS_18_63_port);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => N917, CK => CLK, Q => 
                           n_1640, QN => n1153_port);
   NEXT_REGISTERS_reg_18_62_inst : DLH_X1 port map( G => n12045, D => N3142, Q 
                           => NEXT_REGISTERS_18_62_port);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => N916, CK => CLK, Q => 
                           n_1641, QN => n1154_port);
   NEXT_REGISTERS_reg_18_61_inst : DLH_X1 port map( G => n12045, D => N3141, Q 
                           => NEXT_REGISTERS_18_61_port);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => N915, CK => CLK, Q => 
                           n_1642, QN => n1155_port);
   NEXT_REGISTERS_reg_18_60_inst : DLH_X1 port map( G => n12045, D => N3140, Q 
                           => NEXT_REGISTERS_18_60_port);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => N914, CK => CLK, Q => 
                           n_1643, QN => n1156_port);
   NEXT_REGISTERS_reg_18_59_inst : DLH_X1 port map( G => n12045, D => N3139, Q 
                           => NEXT_REGISTERS_18_59_port);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => N913, CK => CLK, Q => 
                           n_1644, QN => n1157_port);
   NEXT_REGISTERS_reg_18_58_inst : DLH_X1 port map( G => n12045, D => N3138, Q 
                           => NEXT_REGISTERS_18_58_port);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => N912, CK => CLK, Q => 
                           n_1645, QN => n1158_port);
   NEXT_REGISTERS_reg_18_57_inst : DLH_X1 port map( G => n12045, D => N3137, Q 
                           => NEXT_REGISTERS_18_57_port);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => N911, CK => CLK, Q => 
                           n_1646, QN => n1159_port);
   NEXT_REGISTERS_reg_18_56_inst : DLH_X1 port map( G => n12045, D => N3136, Q 
                           => NEXT_REGISTERS_18_56_port);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => N910, CK => CLK, Q => 
                           n_1647, QN => n1160_port);
   NEXT_REGISTERS_reg_18_55_inst : DLH_X1 port map( G => n12045, D => N3135, Q 
                           => NEXT_REGISTERS_18_55_port);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => N909, CK => CLK, Q => 
                           n_1648, QN => n1161_port);
   NEXT_REGISTERS_reg_18_54_inst : DLH_X1 port map( G => n12045, D => N3134, Q 
                           => NEXT_REGISTERS_18_54_port);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => N908, CK => CLK, Q => 
                           n_1649, QN => n1162_port);
   NEXT_REGISTERS_reg_18_53_inst : DLH_X1 port map( G => n12045, D => N3133, Q 
                           => NEXT_REGISTERS_18_53_port);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => N907, CK => CLK, Q => 
                           n_1650, QN => n1163_port);
   NEXT_REGISTERS_reg_18_52_inst : DLH_X1 port map( G => n12046, D => N3132, Q 
                           => NEXT_REGISTERS_18_52_port);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => N906, CK => CLK, Q => 
                           n_1651, QN => n1164_port);
   NEXT_REGISTERS_reg_18_51_inst : DLH_X1 port map( G => n12046, D => N3131, Q 
                           => NEXT_REGISTERS_18_51_port);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => N905, CK => CLK, Q => 
                           n_1652, QN => n1165_port);
   NEXT_REGISTERS_reg_18_50_inst : DLH_X1 port map( G => n12046, D => N3130, Q 
                           => NEXT_REGISTERS_18_50_port);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => N904, CK => CLK, Q => 
                           n_1653, QN => n1166_port);
   NEXT_REGISTERS_reg_18_49_inst : DLH_X1 port map( G => n12046, D => N3129, Q 
                           => NEXT_REGISTERS_18_49_port);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => N903, CK => CLK, Q => 
                           n_1654, QN => n1167_port);
   NEXT_REGISTERS_reg_18_48_inst : DLH_X1 port map( G => n12046, D => N3128, Q 
                           => NEXT_REGISTERS_18_48_port);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => N902, CK => CLK, Q => 
                           n_1655, QN => n1168_port);
   NEXT_REGISTERS_reg_18_47_inst : DLH_X1 port map( G => n12046, D => N3127, Q 
                           => NEXT_REGISTERS_18_47_port);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => N901, CK => CLK, Q => 
                           n_1656, QN => n1169_port);
   NEXT_REGISTERS_reg_18_46_inst : DLH_X1 port map( G => n12046, D => N3126, Q 
                           => NEXT_REGISTERS_18_46_port);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => N900, CK => CLK, Q => 
                           n_1657, QN => n1170_port);
   NEXT_REGISTERS_reg_18_45_inst : DLH_X1 port map( G => n12046, D => N3125, Q 
                           => NEXT_REGISTERS_18_45_port);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => N899, CK => CLK, Q => 
                           n_1658, QN => n1171_port);
   NEXT_REGISTERS_reg_18_44_inst : DLH_X1 port map( G => n12046, D => N3124, Q 
                           => NEXT_REGISTERS_18_44_port);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => N898, CK => CLK, Q => 
                           n_1659, QN => n1172_port);
   NEXT_REGISTERS_reg_18_43_inst : DLH_X1 port map( G => n12046, D => N3123, Q 
                           => NEXT_REGISTERS_18_43_port);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => N897, CK => CLK, Q => 
                           n_1660, QN => n1173_port);
   NEXT_REGISTERS_reg_18_42_inst : DLH_X1 port map( G => n12046, D => N3122, Q 
                           => NEXT_REGISTERS_18_42_port);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => N896, CK => CLK, Q => 
                           n_1661, QN => n1174_port);
   NEXT_REGISTERS_reg_18_41_inst : DLH_X1 port map( G => n12047, D => N3121, Q 
                           => NEXT_REGISTERS_18_41_port);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => N895, CK => CLK, Q => 
                           n_1662, QN => n1175_port);
   NEXT_REGISTERS_reg_18_40_inst : DLH_X1 port map( G => n12047, D => N3120, Q 
                           => NEXT_REGISTERS_18_40_port);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => N894, CK => CLK, Q => 
                           n_1663, QN => n1176_port);
   NEXT_REGISTERS_reg_18_39_inst : DLH_X1 port map( G => n12047, D => N3119, Q 
                           => NEXT_REGISTERS_18_39_port);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => N893, CK => CLK, Q => 
                           n_1664, QN => n1177_port);
   NEXT_REGISTERS_reg_18_38_inst : DLH_X1 port map( G => n12047, D => N3118, Q 
                           => NEXT_REGISTERS_18_38_port);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => N892, CK => CLK, Q => 
                           n_1665, QN => n1178_port);
   NEXT_REGISTERS_reg_18_37_inst : DLH_X1 port map( G => n12047, D => N3117, Q 
                           => NEXT_REGISTERS_18_37_port);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => N891, CK => CLK, Q => 
                           n_1666, QN => n1179_port);
   NEXT_REGISTERS_reg_18_36_inst : DLH_X1 port map( G => n12047, D => N3116, Q 
                           => NEXT_REGISTERS_18_36_port);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => N890, CK => CLK, Q => 
                           n_1667, QN => n1180_port);
   NEXT_REGISTERS_reg_18_35_inst : DLH_X1 port map( G => n12047, D => N3115, Q 
                           => NEXT_REGISTERS_18_35_port);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => N889, CK => CLK, Q => 
                           n_1668, QN => n1181_port);
   NEXT_REGISTERS_reg_18_34_inst : DLH_X1 port map( G => n12047, D => N3114, Q 
                           => NEXT_REGISTERS_18_34_port);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => N888, CK => CLK, Q => 
                           n_1669, QN => n1182_port);
   NEXT_REGISTERS_reg_18_33_inst : DLH_X1 port map( G => n12047, D => N3113, Q 
                           => NEXT_REGISTERS_18_33_port);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => N887, CK => CLK, Q => 
                           n_1670, QN => n1183_port);
   NEXT_REGISTERS_reg_18_32_inst : DLH_X1 port map( G => n12047, D => N3112, Q 
                           => NEXT_REGISTERS_18_32_port);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => N886, CK => CLK, Q => 
                           n_1671, QN => n1184_port);
   NEXT_REGISTERS_reg_18_31_inst : DLH_X1 port map( G => n12047, D => N3111, Q 
                           => NEXT_REGISTERS_18_31_port);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => N885, CK => CLK, Q => 
                           n_1672, QN => n1185_port);
   NEXT_REGISTERS_reg_18_30_inst : DLH_X1 port map( G => n12048, D => N3110, Q 
                           => NEXT_REGISTERS_18_30_port);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => N884, CK => CLK, Q => 
                           n_1673, QN => n1186_port);
   NEXT_REGISTERS_reg_18_29_inst : DLH_X1 port map( G => n12048, D => N3109, Q 
                           => NEXT_REGISTERS_18_29_port);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => N883, CK => CLK, Q => 
                           n_1674, QN => n1187_port);
   NEXT_REGISTERS_reg_18_28_inst : DLH_X1 port map( G => n12048, D => N3108, Q 
                           => NEXT_REGISTERS_18_28_port);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => N882, CK => CLK, Q => 
                           n_1675, QN => n1188_port);
   NEXT_REGISTERS_reg_18_27_inst : DLH_X1 port map( G => n12048, D => N3107, Q 
                           => NEXT_REGISTERS_18_27_port);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => N881, CK => CLK, Q => 
                           n_1676, QN => n1189_port);
   NEXT_REGISTERS_reg_18_26_inst : DLH_X1 port map( G => n12048, D => N3106, Q 
                           => NEXT_REGISTERS_18_26_port);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => N880, CK => CLK, Q => 
                           n_1677, QN => n1190_port);
   NEXT_REGISTERS_reg_18_25_inst : DLH_X1 port map( G => n12048, D => N3105, Q 
                           => NEXT_REGISTERS_18_25_port);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => N879, CK => CLK, Q => 
                           n_1678, QN => n1191_port);
   NEXT_REGISTERS_reg_18_24_inst : DLH_X1 port map( G => n12048, D => N3104, Q 
                           => NEXT_REGISTERS_18_24_port);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => N878, CK => CLK, Q => 
                           n_1679, QN => n1192_port);
   NEXT_REGISTERS_reg_18_23_inst : DLH_X1 port map( G => n12048, D => N3103, Q 
                           => NEXT_REGISTERS_18_23_port);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => N877, CK => CLK, Q => 
                           n_1680, QN => n1193_port);
   NEXT_REGISTERS_reg_18_22_inst : DLH_X1 port map( G => n12048, D => N3102, Q 
                           => NEXT_REGISTERS_18_22_port);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => N876, CK => CLK, Q => 
                           n_1681, QN => n1194_port);
   NEXT_REGISTERS_reg_18_21_inst : DLH_X1 port map( G => n12048, D => N3101, Q 
                           => NEXT_REGISTERS_18_21_port);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => N875, CK => CLK, Q => 
                           n_1682, QN => n1195_port);
   NEXT_REGISTERS_reg_18_20_inst : DLH_X1 port map( G => n12048, D => N3100, Q 
                           => NEXT_REGISTERS_18_20_port);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => N874, CK => CLK, Q => 
                           n_1683, QN => n1196_port);
   NEXT_REGISTERS_reg_18_19_inst : DLH_X1 port map( G => n12049, D => N3099, Q 
                           => NEXT_REGISTERS_18_19_port);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => N873, CK => CLK, Q => 
                           n_1684, QN => n1197_port);
   NEXT_REGISTERS_reg_18_18_inst : DLH_X1 port map( G => n12049, D => N3098, Q 
                           => NEXT_REGISTERS_18_18_port);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => N872, CK => CLK, Q => 
                           n_1685, QN => n1198_port);
   NEXT_REGISTERS_reg_18_17_inst : DLH_X1 port map( G => n12049, D => N3097, Q 
                           => NEXT_REGISTERS_18_17_port);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => N871, CK => CLK, Q => 
                           n_1686, QN => n1199_port);
   NEXT_REGISTERS_reg_18_16_inst : DLH_X1 port map( G => n12049, D => N3096, Q 
                           => NEXT_REGISTERS_18_16_port);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => N870, CK => CLK, Q => 
                           n_1687, QN => n1200_port);
   NEXT_REGISTERS_reg_18_15_inst : DLH_X1 port map( G => n12049, D => N3095, Q 
                           => NEXT_REGISTERS_18_15_port);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => N869, CK => CLK, Q => 
                           n_1688, QN => n1201_port);
   NEXT_REGISTERS_reg_18_14_inst : DLH_X1 port map( G => n12049, D => N3094, Q 
                           => NEXT_REGISTERS_18_14_port);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => N868, CK => CLK, Q => 
                           n_1689, QN => n1202_port);
   NEXT_REGISTERS_reg_18_13_inst : DLH_X1 port map( G => n12049, D => N3093, Q 
                           => NEXT_REGISTERS_18_13_port);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => N867, CK => CLK, Q => 
                           n_1690, QN => n1203_port);
   NEXT_REGISTERS_reg_18_12_inst : DLH_X1 port map( G => n12049, D => N3092, Q 
                           => NEXT_REGISTERS_18_12_port);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => N866, CK => CLK, Q => 
                           n_1691, QN => n1204_port);
   NEXT_REGISTERS_reg_18_11_inst : DLH_X1 port map( G => n12049, D => N3091, Q 
                           => NEXT_REGISTERS_18_11_port);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => N865, CK => CLK, Q => 
                           n_1692, QN => n1205_port);
   NEXT_REGISTERS_reg_18_10_inst : DLH_X1 port map( G => n12049, D => N3090, Q 
                           => NEXT_REGISTERS_18_10_port);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => N864, CK => CLK, Q => 
                           n_1693, QN => n1206_port);
   NEXT_REGISTERS_reg_18_9_inst : DLH_X1 port map( G => n12049, D => N3089, Q 
                           => NEXT_REGISTERS_18_9_port);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => N863, CK => CLK, Q => n_1694
                           , QN => n1207_port);
   NEXT_REGISTERS_reg_18_8_inst : DLH_X1 port map( G => n12050, D => N3088, Q 
                           => NEXT_REGISTERS_18_8_port);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => N862, CK => CLK, Q => n_1695
                           , QN => n1208_port);
   NEXT_REGISTERS_reg_18_7_inst : DLH_X1 port map( G => n12050, D => N3087, Q 
                           => NEXT_REGISTERS_18_7_port);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => N861, CK => CLK, Q => n_1696
                           , QN => n1209_port);
   NEXT_REGISTERS_reg_18_6_inst : DLH_X1 port map( G => n12050, D => N3086, Q 
                           => NEXT_REGISTERS_18_6_port);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => N860, CK => CLK, Q => n_1697
                           , QN => n1210_port);
   NEXT_REGISTERS_reg_18_5_inst : DLH_X1 port map( G => n12050, D => N3085, Q 
                           => NEXT_REGISTERS_18_5_port);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => N859, CK => CLK, Q => n_1698
                           , QN => n1211_port);
   NEXT_REGISTERS_reg_18_4_inst : DLH_X1 port map( G => n12050, D => N3084, Q 
                           => NEXT_REGISTERS_18_4_port);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => N858, CK => CLK, Q => n_1699
                           , QN => n1212_port);
   NEXT_REGISTERS_reg_18_3_inst : DLH_X1 port map( G => n12050, D => N3083, Q 
                           => NEXT_REGISTERS_18_3_port);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => N857, CK => CLK, Q => n_1700
                           , QN => n1213_port);
   NEXT_REGISTERS_reg_18_2_inst : DLH_X1 port map( G => n12050, D => N3082, Q 
                           => NEXT_REGISTERS_18_2_port);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => N856, CK => CLK, Q => n_1701
                           , QN => n1214_port);
   NEXT_REGISTERS_reg_18_1_inst : DLH_X1 port map( G => n12050, D => N3081, Q 
                           => NEXT_REGISTERS_18_1_port);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => N855, CK => CLK, Q => n_1702
                           , QN => n1215_port);
   NEXT_REGISTERS_reg_18_0_inst : DLH_X1 port map( G => n12050, D => N3080, Q 
                           => NEXT_REGISTERS_18_0_port);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => N854, CK => CLK, Q => n_1703
                           , QN => n1216_port);
   NEXT_REGISTERS_reg_19_63_inst : DLH_X1 port map( G => n12054, D => N3078, Q 
                           => NEXT_REGISTERS_19_63_port);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => N853, CK => CLK, Q => 
                           n10286, QN => n1217_port);
   NEXT_REGISTERS_reg_19_62_inst : DLH_X1 port map( G => n12054, D => N3077, Q 
                           => NEXT_REGISTERS_19_62_port);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => N852, CK => CLK, Q => 
                           n10284, QN => n1218_port);
   NEXT_REGISTERS_reg_19_61_inst : DLH_X1 port map( G => n12054, D => N3076, Q 
                           => NEXT_REGISTERS_19_61_port);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => N851, CK => CLK, Q => 
                           n10282, QN => n1219_port);
   NEXT_REGISTERS_reg_19_60_inst : DLH_X1 port map( G => n12054, D => N3075, Q 
                           => NEXT_REGISTERS_19_60_port);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => N850, CK => CLK, Q => 
                           n10280, QN => n1220_port);
   NEXT_REGISTERS_reg_19_59_inst : DLH_X1 port map( G => n12054, D => N3074, Q 
                           => NEXT_REGISTERS_19_59_port);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => N849, CK => CLK, Q => 
                           n10278, QN => n1221_port);
   NEXT_REGISTERS_reg_19_58_inst : DLH_X1 port map( G => n12054, D => N3073, Q 
                           => NEXT_REGISTERS_19_58_port);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => N848, CK => CLK, Q => 
                           n10276, QN => n1222_port);
   NEXT_REGISTERS_reg_19_57_inst : DLH_X1 port map( G => n12054, D => N3072, Q 
                           => NEXT_REGISTERS_19_57_port);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => N847, CK => CLK, Q => 
                           n10274, QN => n1223_port);
   NEXT_REGISTERS_reg_19_56_inst : DLH_X1 port map( G => n12054, D => N3071, Q 
                           => NEXT_REGISTERS_19_56_port);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => N846, CK => CLK, Q => 
                           n10272, QN => n1224_port);
   NEXT_REGISTERS_reg_19_55_inst : DLH_X1 port map( G => n12054, D => N3070, Q 
                           => NEXT_REGISTERS_19_55_port);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => N845, CK => CLK, Q => 
                           n10270, QN => n1225_port);
   NEXT_REGISTERS_reg_19_54_inst : DLH_X1 port map( G => n12054, D => N3069, Q 
                           => NEXT_REGISTERS_19_54_port);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => N844, CK => CLK, Q => 
                           n10268, QN => n1226_port);
   NEXT_REGISTERS_reg_19_53_inst : DLH_X1 port map( G => n12054, D => N3068, Q 
                           => NEXT_REGISTERS_19_53_port);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => N843, CK => CLK, Q => 
                           n10266, QN => n1227_port);
   NEXT_REGISTERS_reg_19_52_inst : DLH_X1 port map( G => n12055, D => N3067, Q 
                           => NEXT_REGISTERS_19_52_port);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => N842, CK => CLK, Q => 
                           n10264, QN => n1228_port);
   NEXT_REGISTERS_reg_19_51_inst : DLH_X1 port map( G => n12055, D => N3066, Q 
                           => NEXT_REGISTERS_19_51_port);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => N841, CK => CLK, Q => 
                           n10262, QN => n1229_port);
   NEXT_REGISTERS_reg_19_50_inst : DLH_X1 port map( G => n12055, D => N3065, Q 
                           => NEXT_REGISTERS_19_50_port);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => N840, CK => CLK, Q => 
                           n10260, QN => n1230_port);
   NEXT_REGISTERS_reg_19_49_inst : DLH_X1 port map( G => n12055, D => N3064, Q 
                           => NEXT_REGISTERS_19_49_port);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => N839, CK => CLK, Q => 
                           n10258, QN => n1231_port);
   NEXT_REGISTERS_reg_19_48_inst : DLH_X1 port map( G => n12055, D => N3063, Q 
                           => NEXT_REGISTERS_19_48_port);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => N838, CK => CLK, Q => 
                           n10256, QN => n1232_port);
   NEXT_REGISTERS_reg_19_47_inst : DLH_X1 port map( G => n12055, D => N3062, Q 
                           => NEXT_REGISTERS_19_47_port);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => N837, CK => CLK, Q => 
                           n10254, QN => n1233_port);
   NEXT_REGISTERS_reg_19_46_inst : DLH_X1 port map( G => n12055, D => N3061, Q 
                           => NEXT_REGISTERS_19_46_port);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => N836, CK => CLK, Q => 
                           n10252, QN => n1234_port);
   NEXT_REGISTERS_reg_19_45_inst : DLH_X1 port map( G => n12055, D => N3060, Q 
                           => NEXT_REGISTERS_19_45_port);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => N835, CK => CLK, Q => 
                           n10250, QN => n1235_port);
   NEXT_REGISTERS_reg_19_44_inst : DLH_X1 port map( G => n12055, D => N3059, Q 
                           => NEXT_REGISTERS_19_44_port);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => N834, CK => CLK, Q => 
                           n10248, QN => n1236_port);
   NEXT_REGISTERS_reg_19_43_inst : DLH_X1 port map( G => n12055, D => N3058, Q 
                           => NEXT_REGISTERS_19_43_port);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => N833, CK => CLK, Q => 
                           n10246, QN => n1237_port);
   NEXT_REGISTERS_reg_19_42_inst : DLH_X1 port map( G => n12055, D => N3057, Q 
                           => NEXT_REGISTERS_19_42_port);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => N832, CK => CLK, Q => 
                           n10244, QN => n1238_port);
   NEXT_REGISTERS_reg_19_41_inst : DLH_X1 port map( G => n12056, D => N3056, Q 
                           => NEXT_REGISTERS_19_41_port);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => N831, CK => CLK, Q => 
                           n10242, QN => n1239_port);
   NEXT_REGISTERS_reg_19_40_inst : DLH_X1 port map( G => n12056, D => N3055, Q 
                           => NEXT_REGISTERS_19_40_port);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => N830, CK => CLK, Q => 
                           n10240, QN => n1240_port);
   NEXT_REGISTERS_reg_19_39_inst : DLH_X1 port map( G => n12056, D => N3054, Q 
                           => NEXT_REGISTERS_19_39_port);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => N829, CK => CLK, Q => 
                           n10238, QN => n1241_port);
   NEXT_REGISTERS_reg_19_38_inst : DLH_X1 port map( G => n12056, D => N3053, Q 
                           => NEXT_REGISTERS_19_38_port);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => N828, CK => CLK, Q => 
                           n10236, QN => n1242_port);
   NEXT_REGISTERS_reg_19_37_inst : DLH_X1 port map( G => n12056, D => N3052, Q 
                           => NEXT_REGISTERS_19_37_port);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => N827, CK => CLK, Q => 
                           n10234, QN => n1243_port);
   NEXT_REGISTERS_reg_19_36_inst : DLH_X1 port map( G => n12056, D => N3051, Q 
                           => NEXT_REGISTERS_19_36_port);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => N826, CK => CLK, Q => 
                           n10232, QN => n1244_port);
   NEXT_REGISTERS_reg_19_35_inst : DLH_X1 port map( G => n12056, D => N3050, Q 
                           => NEXT_REGISTERS_19_35_port);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => N825, CK => CLK, Q => 
                           n10230, QN => n1245_port);
   NEXT_REGISTERS_reg_19_34_inst : DLH_X1 port map( G => n12056, D => N3049, Q 
                           => NEXT_REGISTERS_19_34_port);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => N824, CK => CLK, Q => 
                           n10228, QN => n1246_port);
   NEXT_REGISTERS_reg_19_33_inst : DLH_X1 port map( G => n12056, D => N3048, Q 
                           => NEXT_REGISTERS_19_33_port);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => N823, CK => CLK, Q => 
                           n10226, QN => n1247_port);
   NEXT_REGISTERS_reg_19_32_inst : DLH_X1 port map( G => n12056, D => N3047, Q 
                           => NEXT_REGISTERS_19_32_port);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => N822, CK => CLK, Q => 
                           n10224, QN => n1248_port);
   NEXT_REGISTERS_reg_19_31_inst : DLH_X1 port map( G => n12056, D => N3046, Q 
                           => NEXT_REGISTERS_19_31_port);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => N821, CK => CLK, Q => 
                           n10222, QN => n1249_port);
   NEXT_REGISTERS_reg_19_30_inst : DLH_X1 port map( G => n12057, D => N3045, Q 
                           => NEXT_REGISTERS_19_30_port);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => N820, CK => CLK, Q => 
                           n10220, QN => n1250_port);
   NEXT_REGISTERS_reg_19_29_inst : DLH_X1 port map( G => n12057, D => N3044, Q 
                           => NEXT_REGISTERS_19_29_port);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => N819, CK => CLK, Q => 
                           n10218, QN => n1251_port);
   NEXT_REGISTERS_reg_19_28_inst : DLH_X1 port map( G => n12057, D => N3043, Q 
                           => NEXT_REGISTERS_19_28_port);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => N818, CK => CLK, Q => 
                           n10216, QN => n1252_port);
   NEXT_REGISTERS_reg_19_27_inst : DLH_X1 port map( G => n12057, D => N3042, Q 
                           => NEXT_REGISTERS_19_27_port);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => N817, CK => CLK, Q => 
                           n10214, QN => n1253_port);
   NEXT_REGISTERS_reg_19_26_inst : DLH_X1 port map( G => n12057, D => N3041, Q 
                           => NEXT_REGISTERS_19_26_port);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => N816, CK => CLK, Q => 
                           n10212, QN => n1254_port);
   NEXT_REGISTERS_reg_19_25_inst : DLH_X1 port map( G => n12057, D => N3040, Q 
                           => NEXT_REGISTERS_19_25_port);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => N815, CK => CLK, Q => 
                           n10210, QN => n1255_port);
   NEXT_REGISTERS_reg_19_24_inst : DLH_X1 port map( G => n12057, D => N3039, Q 
                           => NEXT_REGISTERS_19_24_port);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => N814, CK => CLK, Q => 
                           n10208, QN => n1256_port);
   NEXT_REGISTERS_reg_19_23_inst : DLH_X1 port map( G => n12057, D => N3038, Q 
                           => NEXT_REGISTERS_19_23_port);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => N813, CK => CLK, Q => 
                           n10206, QN => n1257_port);
   NEXT_REGISTERS_reg_19_22_inst : DLH_X1 port map( G => n12057, D => N3037, Q 
                           => NEXT_REGISTERS_19_22_port);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => N812, CK => CLK, Q => 
                           n10204, QN => n1258_port);
   NEXT_REGISTERS_reg_19_21_inst : DLH_X1 port map( G => n12057, D => N3036, Q 
                           => NEXT_REGISTERS_19_21_port);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => N811, CK => CLK, Q => 
                           n10202, QN => n1259_port);
   NEXT_REGISTERS_reg_19_20_inst : DLH_X1 port map( G => n12057, D => N3035, Q 
                           => NEXT_REGISTERS_19_20_port);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => N810, CK => CLK, Q => 
                           n10200, QN => n1260_port);
   NEXT_REGISTERS_reg_19_19_inst : DLH_X1 port map( G => n12058, D => N3034, Q 
                           => NEXT_REGISTERS_19_19_port);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => N809, CK => CLK, Q => 
                           n10198, QN => n1261_port);
   NEXT_REGISTERS_reg_19_18_inst : DLH_X1 port map( G => n12058, D => N3033, Q 
                           => NEXT_REGISTERS_19_18_port);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => N808, CK => CLK, Q => 
                           n10196, QN => n1262_port);
   NEXT_REGISTERS_reg_19_17_inst : DLH_X1 port map( G => n12058, D => N3032, Q 
                           => NEXT_REGISTERS_19_17_port);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => N807, CK => CLK, Q => 
                           n10194, QN => n1263_port);
   NEXT_REGISTERS_reg_19_16_inst : DLH_X1 port map( G => n12058, D => N3031, Q 
                           => NEXT_REGISTERS_19_16_port);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => N806, CK => CLK, Q => 
                           n10192, QN => n1264_port);
   NEXT_REGISTERS_reg_19_15_inst : DLH_X1 port map( G => n12058, D => N3030, Q 
                           => NEXT_REGISTERS_19_15_port);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => N805, CK => CLK, Q => 
                           n10190, QN => n1265_port);
   NEXT_REGISTERS_reg_19_14_inst : DLH_X1 port map( G => n12058, D => N3029, Q 
                           => NEXT_REGISTERS_19_14_port);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => N804, CK => CLK, Q => 
                           n10188, QN => n1266_port);
   NEXT_REGISTERS_reg_19_13_inst : DLH_X1 port map( G => n12058, D => N3028, Q 
                           => NEXT_REGISTERS_19_13_port);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => N803, CK => CLK, Q => 
                           n10186, QN => n1267_port);
   NEXT_REGISTERS_reg_19_12_inst : DLH_X1 port map( G => n12058, D => N3027, Q 
                           => NEXT_REGISTERS_19_12_port);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => N802, CK => CLK, Q => 
                           n10184, QN => n1268_port);
   NEXT_REGISTERS_reg_19_11_inst : DLH_X1 port map( G => n12058, D => N3026, Q 
                           => NEXT_REGISTERS_19_11_port);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => N801, CK => CLK, Q => 
                           n10182, QN => n1269_port);
   NEXT_REGISTERS_reg_19_10_inst : DLH_X1 port map( G => n12058, D => N3025, Q 
                           => NEXT_REGISTERS_19_10_port);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => N800, CK => CLK, Q => 
                           n10180, QN => n1270_port);
   NEXT_REGISTERS_reg_19_9_inst : DLH_X1 port map( G => n12058, D => N3024, Q 
                           => NEXT_REGISTERS_19_9_port);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => N799, CK => CLK, Q => n10178
                           , QN => n1271_port);
   NEXT_REGISTERS_reg_19_8_inst : DLH_X1 port map( G => n12059, D => N3023, Q 
                           => NEXT_REGISTERS_19_8_port);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => N798, CK => CLK, Q => n10176
                           , QN => n1272_port);
   NEXT_REGISTERS_reg_19_7_inst : DLH_X1 port map( G => n12059, D => N3022, Q 
                           => NEXT_REGISTERS_19_7_port);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => N797, CK => CLK, Q => n10174
                           , QN => n1273_port);
   NEXT_REGISTERS_reg_19_6_inst : DLH_X1 port map( G => n12059, D => N3021, Q 
                           => NEXT_REGISTERS_19_6_port);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => N796, CK => CLK, Q => n10172
                           , QN => n1274_port);
   NEXT_REGISTERS_reg_19_5_inst : DLH_X1 port map( G => n12059, D => N3020, Q 
                           => NEXT_REGISTERS_19_5_port);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => N795, CK => CLK, Q => n10170
                           , QN => n1275_port);
   NEXT_REGISTERS_reg_19_4_inst : DLH_X1 port map( G => n12059, D => N3019, Q 
                           => NEXT_REGISTERS_19_4_port);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => N794, CK => CLK, Q => n10168
                           , QN => n1276_port);
   NEXT_REGISTERS_reg_19_3_inst : DLH_X1 port map( G => n12059, D => N3018, Q 
                           => NEXT_REGISTERS_19_3_port);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => N793, CK => CLK, Q => n10166
                           , QN => n1277_port);
   NEXT_REGISTERS_reg_19_2_inst : DLH_X1 port map( G => n12059, D => N3017, Q 
                           => NEXT_REGISTERS_19_2_port);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => N792, CK => CLK, Q => n10164
                           , QN => n1278_port);
   NEXT_REGISTERS_reg_19_1_inst : DLH_X1 port map( G => n12059, D => N3016, Q 
                           => NEXT_REGISTERS_19_1_port);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => N791, CK => CLK, Q => n10162
                           , QN => n1279_port);
   NEXT_REGISTERS_reg_19_0_inst : DLH_X1 port map( G => n12059, D => N3015, Q 
                           => NEXT_REGISTERS_19_0_port);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => N790, CK => CLK, Q => n10160
                           , QN => n1280_port);
   NEXT_REGISTERS_reg_20_63_inst : DLH_X1 port map( G => n12063, D => N3013, Q 
                           => NEXT_REGISTERS_20_63_port);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => N789, CK => CLK, Q => n9838
                           , QN => n1281_port);
   NEXT_REGISTERS_reg_20_62_inst : DLH_X1 port map( G => n12063, D => N3012, Q 
                           => NEXT_REGISTERS_20_62_port);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => N788, CK => CLK, Q => n9836
                           , QN => n1282_port);
   NEXT_REGISTERS_reg_20_61_inst : DLH_X1 port map( G => n12063, D => N3011, Q 
                           => NEXT_REGISTERS_20_61_port);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => N787, CK => CLK, Q => n9834
                           , QN => n1283_port);
   NEXT_REGISTERS_reg_20_60_inst : DLH_X1 port map( G => n12063, D => N3010, Q 
                           => NEXT_REGISTERS_20_60_port);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => N786, CK => CLK, Q => n9832
                           , QN => n1284_port);
   NEXT_REGISTERS_reg_20_59_inst : DLH_X1 port map( G => n12063, D => N3009, Q 
                           => NEXT_REGISTERS_20_59_port);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => N785, CK => CLK, Q => n9830
                           , QN => n1285_port);
   NEXT_REGISTERS_reg_20_58_inst : DLH_X1 port map( G => n12063, D => N3008, Q 
                           => NEXT_REGISTERS_20_58_port);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => N784, CK => CLK, Q => n9828
                           , QN => n1286_port);
   NEXT_REGISTERS_reg_20_57_inst : DLH_X1 port map( G => n12063, D => N3007, Q 
                           => NEXT_REGISTERS_20_57_port);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => N783, CK => CLK, Q => n9826
                           , QN => n1287_port);
   NEXT_REGISTERS_reg_20_56_inst : DLH_X1 port map( G => n12063, D => N3006, Q 
                           => NEXT_REGISTERS_20_56_port);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => N782, CK => CLK, Q => n9824
                           , QN => n1288_port);
   NEXT_REGISTERS_reg_20_55_inst : DLH_X1 port map( G => n12063, D => N3005, Q 
                           => NEXT_REGISTERS_20_55_port);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => N781, CK => CLK, Q => n9822
                           , QN => n1289_port);
   NEXT_REGISTERS_reg_20_54_inst : DLH_X1 port map( G => n12063, D => N3004, Q 
                           => NEXT_REGISTERS_20_54_port);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => N780, CK => CLK, Q => n9820
                           , QN => n1290_port);
   NEXT_REGISTERS_reg_20_53_inst : DLH_X1 port map( G => n12063, D => N3003, Q 
                           => NEXT_REGISTERS_20_53_port);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => N779, CK => CLK, Q => n9818
                           , QN => n1291_port);
   NEXT_REGISTERS_reg_20_52_inst : DLH_X1 port map( G => n12064, D => N3002, Q 
                           => NEXT_REGISTERS_20_52_port);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => N778, CK => CLK, Q => n9816
                           , QN => n1292_port);
   NEXT_REGISTERS_reg_20_51_inst : DLH_X1 port map( G => n12064, D => N3001, Q 
                           => NEXT_REGISTERS_20_51_port);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => N777, CK => CLK, Q => n9814
                           , QN => n1293_port);
   NEXT_REGISTERS_reg_20_50_inst : DLH_X1 port map( G => n12064, D => N3000, Q 
                           => NEXT_REGISTERS_20_50_port);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => N776, CK => CLK, Q => n9812
                           , QN => n1294_port);
   NEXT_REGISTERS_reg_20_49_inst : DLH_X1 port map( G => n12064, D => N2999, Q 
                           => NEXT_REGISTERS_20_49_port);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => N775, CK => CLK, Q => n9810
                           , QN => n1295_port);
   NEXT_REGISTERS_reg_20_48_inst : DLH_X1 port map( G => n12064, D => N2998, Q 
                           => NEXT_REGISTERS_20_48_port);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => N774, CK => CLK, Q => n9808
                           , QN => n1296_port);
   NEXT_REGISTERS_reg_20_47_inst : DLH_X1 port map( G => n12064, D => N2997, Q 
                           => NEXT_REGISTERS_20_47_port);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => N773, CK => CLK, Q => n9806
                           , QN => n1297_port);
   NEXT_REGISTERS_reg_20_46_inst : DLH_X1 port map( G => n12064, D => N2996, Q 
                           => NEXT_REGISTERS_20_46_port);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => N772, CK => CLK, Q => n9804
                           , QN => n1298_port);
   NEXT_REGISTERS_reg_20_45_inst : DLH_X1 port map( G => n12064, D => N2995, Q 
                           => NEXT_REGISTERS_20_45_port);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => N771, CK => CLK, Q => n9802
                           , QN => n1299_port);
   NEXT_REGISTERS_reg_20_44_inst : DLH_X1 port map( G => n12064, D => N2994, Q 
                           => NEXT_REGISTERS_20_44_port);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => N770, CK => CLK, Q => n9800
                           , QN => n1300_port);
   NEXT_REGISTERS_reg_20_43_inst : DLH_X1 port map( G => n12064, D => N2993, Q 
                           => NEXT_REGISTERS_20_43_port);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => N769, CK => CLK, Q => n9798
                           , QN => n1301_port);
   NEXT_REGISTERS_reg_20_42_inst : DLH_X1 port map( G => n12064, D => N2992, Q 
                           => NEXT_REGISTERS_20_42_port);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => N768, CK => CLK, Q => n9796
                           , QN => n1302_port);
   NEXT_REGISTERS_reg_20_41_inst : DLH_X1 port map( G => n12065, D => N2991, Q 
                           => NEXT_REGISTERS_20_41_port);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => N767, CK => CLK, Q => n9794
                           , QN => n1303_port);
   NEXT_REGISTERS_reg_20_40_inst : DLH_X1 port map( G => n12065, D => N2990, Q 
                           => NEXT_REGISTERS_20_40_port);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => N766, CK => CLK, Q => n9792
                           , QN => n1304_port);
   NEXT_REGISTERS_reg_20_39_inst : DLH_X1 port map( G => n12065, D => N2989, Q 
                           => NEXT_REGISTERS_20_39_port);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => N765, CK => CLK, Q => n9790
                           , QN => n1305_port);
   NEXT_REGISTERS_reg_20_38_inst : DLH_X1 port map( G => n12065, D => N2988, Q 
                           => NEXT_REGISTERS_20_38_port);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => N764, CK => CLK, Q => n9788
                           , QN => n1306_port);
   NEXT_REGISTERS_reg_20_37_inst : DLH_X1 port map( G => n12065, D => N2987, Q 
                           => NEXT_REGISTERS_20_37_port);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => N763, CK => CLK, Q => n9786
                           , QN => n1307_port);
   NEXT_REGISTERS_reg_20_36_inst : DLH_X1 port map( G => n12065, D => N2986, Q 
                           => NEXT_REGISTERS_20_36_port);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => N762, CK => CLK, Q => n9784
                           , QN => n1308_port);
   NEXT_REGISTERS_reg_20_35_inst : DLH_X1 port map( G => n12065, D => N2985, Q 
                           => NEXT_REGISTERS_20_35_port);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => N761, CK => CLK, Q => n9782
                           , QN => n1309_port);
   NEXT_REGISTERS_reg_20_34_inst : DLH_X1 port map( G => n12065, D => N2984, Q 
                           => NEXT_REGISTERS_20_34_port);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => N760, CK => CLK, Q => n9780
                           , QN => n1310_port);
   NEXT_REGISTERS_reg_20_33_inst : DLH_X1 port map( G => n12065, D => N2983, Q 
                           => NEXT_REGISTERS_20_33_port);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => N759, CK => CLK, Q => n9778
                           , QN => n1311_port);
   NEXT_REGISTERS_reg_20_32_inst : DLH_X1 port map( G => n12065, D => N2982, Q 
                           => NEXT_REGISTERS_20_32_port);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => N758, CK => CLK, Q => n9776
                           , QN => n1312_port);
   NEXT_REGISTERS_reg_20_31_inst : DLH_X1 port map( G => n12065, D => N2981, Q 
                           => NEXT_REGISTERS_20_31_port);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => N757, CK => CLK, Q => n9774
                           , QN => n1313_port);
   NEXT_REGISTERS_reg_20_30_inst : DLH_X1 port map( G => n12066, D => N2980, Q 
                           => NEXT_REGISTERS_20_30_port);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => N756, CK => CLK, Q => n9772
                           , QN => n1314_port);
   NEXT_REGISTERS_reg_20_29_inst : DLH_X1 port map( G => n12066, D => N2979, Q 
                           => NEXT_REGISTERS_20_29_port);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => N755, CK => CLK, Q => n9770
                           , QN => n1315_port);
   NEXT_REGISTERS_reg_20_28_inst : DLH_X1 port map( G => n12066, D => N2978, Q 
                           => NEXT_REGISTERS_20_28_port);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => N754, CK => CLK, Q => n9768
                           , QN => n1316_port);
   NEXT_REGISTERS_reg_20_27_inst : DLH_X1 port map( G => n12066, D => N2977, Q 
                           => NEXT_REGISTERS_20_27_port);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => N753, CK => CLK, Q => n9766
                           , QN => n1317_port);
   NEXT_REGISTERS_reg_20_26_inst : DLH_X1 port map( G => n12066, D => N2976, Q 
                           => NEXT_REGISTERS_20_26_port);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => N752, CK => CLK, Q => n9764
                           , QN => n1318_port);
   NEXT_REGISTERS_reg_20_25_inst : DLH_X1 port map( G => n12066, D => N2975, Q 
                           => NEXT_REGISTERS_20_25_port);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => N751, CK => CLK, Q => n9762
                           , QN => n1319_port);
   NEXT_REGISTERS_reg_20_24_inst : DLH_X1 port map( G => n12066, D => N2974, Q 
                           => NEXT_REGISTERS_20_24_port);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => N750, CK => CLK, Q => n9760
                           , QN => n1320_port);
   NEXT_REGISTERS_reg_20_23_inst : DLH_X1 port map( G => n12066, D => N2973, Q 
                           => NEXT_REGISTERS_20_23_port);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => N749, CK => CLK, Q => n9758
                           , QN => n1321_port);
   NEXT_REGISTERS_reg_20_22_inst : DLH_X1 port map( G => n12066, D => N2972, Q 
                           => NEXT_REGISTERS_20_22_port);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => N748, CK => CLK, Q => n9756
                           , QN => n1322_port);
   NEXT_REGISTERS_reg_20_21_inst : DLH_X1 port map( G => n12066, D => N2971, Q 
                           => NEXT_REGISTERS_20_21_port);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => N747, CK => CLK, Q => n9754
                           , QN => n1323_port);
   NEXT_REGISTERS_reg_20_20_inst : DLH_X1 port map( G => n12066, D => N2970, Q 
                           => NEXT_REGISTERS_20_20_port);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => N746, CK => CLK, Q => n9752
                           , QN => n1324_port);
   NEXT_REGISTERS_reg_20_19_inst : DLH_X1 port map( G => n12067, D => N2969, Q 
                           => NEXT_REGISTERS_20_19_port);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => N745, CK => CLK, Q => n9750
                           , QN => n1325_port);
   NEXT_REGISTERS_reg_20_18_inst : DLH_X1 port map( G => n12067, D => N2968, Q 
                           => NEXT_REGISTERS_20_18_port);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => N744, CK => CLK, Q => n9748
                           , QN => n1326_port);
   NEXT_REGISTERS_reg_20_17_inst : DLH_X1 port map( G => n12067, D => N2967, Q 
                           => NEXT_REGISTERS_20_17_port);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => N743, CK => CLK, Q => n9746
                           , QN => n1327_port);
   NEXT_REGISTERS_reg_20_16_inst : DLH_X1 port map( G => n12067, D => N2966, Q 
                           => NEXT_REGISTERS_20_16_port);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => N742, CK => CLK, Q => n9744
                           , QN => n1328_port);
   NEXT_REGISTERS_reg_20_15_inst : DLH_X1 port map( G => n12067, D => N2965, Q 
                           => NEXT_REGISTERS_20_15_port);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => N741, CK => CLK, Q => n9742
                           , QN => n1329_port);
   NEXT_REGISTERS_reg_20_14_inst : DLH_X1 port map( G => n12067, D => N2964, Q 
                           => NEXT_REGISTERS_20_14_port);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => N740, CK => CLK, Q => n9740
                           , QN => n1330_port);
   NEXT_REGISTERS_reg_20_13_inst : DLH_X1 port map( G => n12067, D => N2963, Q 
                           => NEXT_REGISTERS_20_13_port);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => N739, CK => CLK, Q => n9738
                           , QN => n1331_port);
   NEXT_REGISTERS_reg_20_12_inst : DLH_X1 port map( G => n12067, D => N2962, Q 
                           => NEXT_REGISTERS_20_12_port);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => N738, CK => CLK, Q => n9736
                           , QN => n1332_port);
   NEXT_REGISTERS_reg_20_11_inst : DLH_X1 port map( G => n12067, D => N2961, Q 
                           => NEXT_REGISTERS_20_11_port);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => N737, CK => CLK, Q => n9734
                           , QN => n1333_port);
   NEXT_REGISTERS_reg_20_10_inst : DLH_X1 port map( G => n12067, D => N2960, Q 
                           => NEXT_REGISTERS_20_10_port);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => N736, CK => CLK, Q => n9732
                           , QN => n1334_port);
   NEXT_REGISTERS_reg_20_9_inst : DLH_X1 port map( G => n12067, D => N2959, Q 
                           => NEXT_REGISTERS_20_9_port);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => N735, CK => CLK, Q => n9730,
                           QN => n1335_port);
   NEXT_REGISTERS_reg_20_8_inst : DLH_X1 port map( G => n12068, D => N2958, Q 
                           => NEXT_REGISTERS_20_8_port);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => N734, CK => CLK, Q => n9728,
                           QN => n1336_port);
   NEXT_REGISTERS_reg_20_7_inst : DLH_X1 port map( G => n12068, D => N2957, Q 
                           => NEXT_REGISTERS_20_7_port);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => N733, CK => CLK, Q => n9726,
                           QN => n1337_port);
   NEXT_REGISTERS_reg_20_6_inst : DLH_X1 port map( G => n12068, D => N2956, Q 
                           => NEXT_REGISTERS_20_6_port);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => N732, CK => CLK, Q => n9724,
                           QN => n1338_port);
   NEXT_REGISTERS_reg_20_5_inst : DLH_X1 port map( G => n12068, D => N2955, Q 
                           => NEXT_REGISTERS_20_5_port);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => N731, CK => CLK, Q => n9722,
                           QN => n1339_port);
   NEXT_REGISTERS_reg_20_4_inst : DLH_X1 port map( G => n12068, D => N2954, Q 
                           => NEXT_REGISTERS_20_4_port);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => N730, CK => CLK, Q => n9720,
                           QN => n1340_port);
   NEXT_REGISTERS_reg_20_3_inst : DLH_X1 port map( G => n12068, D => N2953, Q 
                           => NEXT_REGISTERS_20_3_port);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => N729, CK => CLK, Q => n9718,
                           QN => n1341_port);
   NEXT_REGISTERS_reg_20_2_inst : DLH_X1 port map( G => n12068, D => N2952, Q 
                           => NEXT_REGISTERS_20_2_port);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => N728, CK => CLK, Q => n9716,
                           QN => n1342_port);
   NEXT_REGISTERS_reg_20_1_inst : DLH_X1 port map( G => n12068, D => N2951, Q 
                           => NEXT_REGISTERS_20_1_port);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => N727, CK => CLK, Q => n9714,
                           QN => n1343_port);
   NEXT_REGISTERS_reg_20_0_inst : DLH_X1 port map( G => n12068, D => N2950, Q 
                           => NEXT_REGISTERS_20_0_port);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => N726, CK => CLK, Q => n9712,
                           QN => n1344_port);
   NEXT_REGISTERS_reg_21_63_inst : DLH_X1 port map( G => n12072, D => N2948, Q 
                           => NEXT_REGISTERS_21_63_port);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => N725, CK => CLK, Q => 
                           n_1704, QN => n1345_port);
   NEXT_REGISTERS_reg_21_62_inst : DLH_X1 port map( G => n12072, D => N2947, Q 
                           => NEXT_REGISTERS_21_62_port);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => N724, CK => CLK, Q => 
                           n_1705, QN => n1346_port);
   NEXT_REGISTERS_reg_21_61_inst : DLH_X1 port map( G => n12072, D => N2946, Q 
                           => NEXT_REGISTERS_21_61_port);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => N723, CK => CLK, Q => 
                           n_1706, QN => n1347_port);
   NEXT_REGISTERS_reg_21_60_inst : DLH_X1 port map( G => n12072, D => N2945, Q 
                           => NEXT_REGISTERS_21_60_port);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => N722, CK => CLK, Q => 
                           n_1707, QN => n1348_port);
   NEXT_REGISTERS_reg_21_59_inst : DLH_X1 port map( G => n12072, D => N2944, Q 
                           => NEXT_REGISTERS_21_59_port);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => N721, CK => CLK, Q => 
                           n_1708, QN => n1349_port);
   NEXT_REGISTERS_reg_21_58_inst : DLH_X1 port map( G => n12072, D => N2943, Q 
                           => NEXT_REGISTERS_21_58_port);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => N720, CK => CLK, Q => 
                           n_1709, QN => n1350_port);
   NEXT_REGISTERS_reg_21_57_inst : DLH_X1 port map( G => n12072, D => N2942, Q 
                           => NEXT_REGISTERS_21_57_port);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => N719, CK => CLK, Q => 
                           n_1710, QN => n1351_port);
   NEXT_REGISTERS_reg_21_56_inst : DLH_X1 port map( G => n12072, D => N2941, Q 
                           => NEXT_REGISTERS_21_56_port);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => N718, CK => CLK, Q => 
                           n_1711, QN => n1352_port);
   NEXT_REGISTERS_reg_21_55_inst : DLH_X1 port map( G => n12072, D => N2940, Q 
                           => NEXT_REGISTERS_21_55_port);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => N717, CK => CLK, Q => 
                           n_1712, QN => n1353_port);
   NEXT_REGISTERS_reg_21_54_inst : DLH_X1 port map( G => n12072, D => N2939, Q 
                           => NEXT_REGISTERS_21_54_port);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => N716, CK => CLK, Q => 
                           n_1713, QN => n1354_port);
   NEXT_REGISTERS_reg_21_53_inst : DLH_X1 port map( G => n12072, D => N2938, Q 
                           => NEXT_REGISTERS_21_53_port);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => N715, CK => CLK, Q => 
                           n_1714, QN => n1355_port);
   NEXT_REGISTERS_reg_21_52_inst : DLH_X1 port map( G => n12073, D => N2937, Q 
                           => NEXT_REGISTERS_21_52_port);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => N714, CK => CLK, Q => 
                           n_1715, QN => n1356_port);
   NEXT_REGISTERS_reg_21_51_inst : DLH_X1 port map( G => n12073, D => N2936, Q 
                           => NEXT_REGISTERS_21_51_port);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => N713, CK => CLK, Q => 
                           n_1716, QN => n1357_port);
   NEXT_REGISTERS_reg_21_50_inst : DLH_X1 port map( G => n12073, D => N2935, Q 
                           => NEXT_REGISTERS_21_50_port);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => N712, CK => CLK, Q => 
                           n_1717, QN => n1358_port);
   NEXT_REGISTERS_reg_21_49_inst : DLH_X1 port map( G => n12073, D => N2934, Q 
                           => NEXT_REGISTERS_21_49_port);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => N711, CK => CLK, Q => 
                           n_1718, QN => n1359_port);
   NEXT_REGISTERS_reg_21_48_inst : DLH_X1 port map( G => n12073, D => N2933, Q 
                           => NEXT_REGISTERS_21_48_port);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => N710, CK => CLK, Q => 
                           n_1719, QN => n1360_port);
   NEXT_REGISTERS_reg_21_47_inst : DLH_X1 port map( G => n12073, D => N2932, Q 
                           => NEXT_REGISTERS_21_47_port);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => N709, CK => CLK, Q => 
                           n_1720, QN => n1361_port);
   NEXT_REGISTERS_reg_21_46_inst : DLH_X1 port map( G => n12073, D => N2931, Q 
                           => NEXT_REGISTERS_21_46_port);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => N708, CK => CLK, Q => 
                           n_1721, QN => n1362_port);
   NEXT_REGISTERS_reg_21_45_inst : DLH_X1 port map( G => n12073, D => N2930, Q 
                           => NEXT_REGISTERS_21_45_port);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => N707, CK => CLK, Q => 
                           n_1722, QN => n1363_port);
   NEXT_REGISTERS_reg_21_44_inst : DLH_X1 port map( G => n12073, D => N2929, Q 
                           => NEXT_REGISTERS_21_44_port);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => N706, CK => CLK, Q => 
                           n_1723, QN => n1364_port);
   NEXT_REGISTERS_reg_21_43_inst : DLH_X1 port map( G => n12073, D => N2928, Q 
                           => NEXT_REGISTERS_21_43_port);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => N705, CK => CLK, Q => 
                           n_1724, QN => n1365_port);
   NEXT_REGISTERS_reg_21_42_inst : DLH_X1 port map( G => n12073, D => N2927, Q 
                           => NEXT_REGISTERS_21_42_port);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => N704, CK => CLK, Q => 
                           n_1725, QN => n1366_port);
   NEXT_REGISTERS_reg_21_41_inst : DLH_X1 port map( G => n12074, D => N2926, Q 
                           => NEXT_REGISTERS_21_41_port);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => N703, CK => CLK, Q => 
                           n_1726, QN => n1367_port);
   NEXT_REGISTERS_reg_21_40_inst : DLH_X1 port map( G => n12074, D => N2925, Q 
                           => NEXT_REGISTERS_21_40_port);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => N702, CK => CLK, Q => 
                           n_1727, QN => n1368_port);
   NEXT_REGISTERS_reg_21_39_inst : DLH_X1 port map( G => n12074, D => N2924, Q 
                           => NEXT_REGISTERS_21_39_port);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => N701, CK => CLK, Q => 
                           n_1728, QN => n1369_port);
   NEXT_REGISTERS_reg_21_38_inst : DLH_X1 port map( G => n12074, D => N2923, Q 
                           => NEXT_REGISTERS_21_38_port);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => N700, CK => CLK, Q => 
                           n_1729, QN => n1370_port);
   NEXT_REGISTERS_reg_21_37_inst : DLH_X1 port map( G => n12074, D => N2922, Q 
                           => NEXT_REGISTERS_21_37_port);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => N699, CK => CLK, Q => 
                           n_1730, QN => n1371_port);
   NEXT_REGISTERS_reg_21_36_inst : DLH_X1 port map( G => n12074, D => N2921, Q 
                           => NEXT_REGISTERS_21_36_port);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => N698, CK => CLK, Q => 
                           n_1731, QN => n1372_port);
   NEXT_REGISTERS_reg_21_35_inst : DLH_X1 port map( G => n12074, D => N2920, Q 
                           => NEXT_REGISTERS_21_35_port);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => N697, CK => CLK, Q => 
                           n_1732, QN => n1373_port);
   NEXT_REGISTERS_reg_21_34_inst : DLH_X1 port map( G => n12074, D => N2919, Q 
                           => NEXT_REGISTERS_21_34_port);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => N696, CK => CLK, Q => 
                           n_1733, QN => n1374_port);
   NEXT_REGISTERS_reg_21_33_inst : DLH_X1 port map( G => n12074, D => N2918, Q 
                           => NEXT_REGISTERS_21_33_port);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => N695, CK => CLK, Q => 
                           n_1734, QN => n1375_port);
   NEXT_REGISTERS_reg_21_32_inst : DLH_X1 port map( G => n12074, D => N2917, Q 
                           => NEXT_REGISTERS_21_32_port);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => N694, CK => CLK, Q => 
                           n_1735, QN => n1376_port);
   NEXT_REGISTERS_reg_21_31_inst : DLH_X1 port map( G => n12074, D => N2916, Q 
                           => NEXT_REGISTERS_21_31_port);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => N693, CK => CLK, Q => 
                           n_1736, QN => n1377_port);
   NEXT_REGISTERS_reg_21_30_inst : DLH_X1 port map( G => n12075, D => N2915, Q 
                           => NEXT_REGISTERS_21_30_port);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => N692, CK => CLK, Q => 
                           n_1737, QN => n1378_port);
   NEXT_REGISTERS_reg_21_29_inst : DLH_X1 port map( G => n12075, D => N2914, Q 
                           => NEXT_REGISTERS_21_29_port);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => N691, CK => CLK, Q => 
                           n_1738, QN => n1379_port);
   NEXT_REGISTERS_reg_21_28_inst : DLH_X1 port map( G => n12075, D => N2913, Q 
                           => NEXT_REGISTERS_21_28_port);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => N690, CK => CLK, Q => 
                           n_1739, QN => n1380_port);
   NEXT_REGISTERS_reg_21_27_inst : DLH_X1 port map( G => n12075, D => N2912, Q 
                           => NEXT_REGISTERS_21_27_port);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => N689, CK => CLK, Q => 
                           n_1740, QN => n1381_port);
   NEXT_REGISTERS_reg_21_26_inst : DLH_X1 port map( G => n12075, D => N2911, Q 
                           => NEXT_REGISTERS_21_26_port);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => N688, CK => CLK, Q => 
                           n_1741, QN => n1382_port);
   NEXT_REGISTERS_reg_21_25_inst : DLH_X1 port map( G => n12075, D => N2910, Q 
                           => NEXT_REGISTERS_21_25_port);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => N687, CK => CLK, Q => 
                           n_1742, QN => n1383_port);
   NEXT_REGISTERS_reg_21_24_inst : DLH_X1 port map( G => n12075, D => N2909, Q 
                           => NEXT_REGISTERS_21_24_port);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => N686, CK => CLK, Q => 
                           n_1743, QN => n1384_port);
   NEXT_REGISTERS_reg_21_23_inst : DLH_X1 port map( G => n12075, D => N2908, Q 
                           => NEXT_REGISTERS_21_23_port);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => N685, CK => CLK, Q => 
                           n_1744, QN => n1385_port);
   NEXT_REGISTERS_reg_21_22_inst : DLH_X1 port map( G => n12075, D => N2907, Q 
                           => NEXT_REGISTERS_21_22_port);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => N684, CK => CLK, Q => 
                           n_1745, QN => n1386_port);
   NEXT_REGISTERS_reg_21_21_inst : DLH_X1 port map( G => n12075, D => N2906, Q 
                           => NEXT_REGISTERS_21_21_port);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => N683, CK => CLK, Q => 
                           n_1746, QN => n1387_port);
   NEXT_REGISTERS_reg_21_20_inst : DLH_X1 port map( G => n12075, D => N2905, Q 
                           => NEXT_REGISTERS_21_20_port);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => N682, CK => CLK, Q => 
                           n_1747, QN => n1388_port);
   NEXT_REGISTERS_reg_21_19_inst : DLH_X1 port map( G => n12076, D => N2904, Q 
                           => NEXT_REGISTERS_21_19_port);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => N681, CK => CLK, Q => 
                           n_1748, QN => n1389_port);
   NEXT_REGISTERS_reg_21_18_inst : DLH_X1 port map( G => n12076, D => N2903, Q 
                           => NEXT_REGISTERS_21_18_port);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => N680, CK => CLK, Q => 
                           n_1749, QN => n1390_port);
   NEXT_REGISTERS_reg_21_17_inst : DLH_X1 port map( G => n12076, D => N2902, Q 
                           => NEXT_REGISTERS_21_17_port);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => N679, CK => CLK, Q => 
                           n_1750, QN => n1391_port);
   NEXT_REGISTERS_reg_21_16_inst : DLH_X1 port map( G => n12076, D => N2901, Q 
                           => NEXT_REGISTERS_21_16_port);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => N678, CK => CLK, Q => 
                           n_1751, QN => n1392_port);
   NEXT_REGISTERS_reg_21_15_inst : DLH_X1 port map( G => n12076, D => N2900, Q 
                           => NEXT_REGISTERS_21_15_port);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => N677, CK => CLK, Q => 
                           n_1752, QN => n1393_port);
   NEXT_REGISTERS_reg_21_14_inst : DLH_X1 port map( G => n12076, D => N2899, Q 
                           => NEXT_REGISTERS_21_14_port);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => N676, CK => CLK, Q => 
                           n_1753, QN => n1394_port);
   NEXT_REGISTERS_reg_21_13_inst : DLH_X1 port map( G => n12076, D => N2898, Q 
                           => NEXT_REGISTERS_21_13_port);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => N675, CK => CLK, Q => 
                           n_1754, QN => n1395_port);
   NEXT_REGISTERS_reg_21_12_inst : DLH_X1 port map( G => n12076, D => N2897, Q 
                           => NEXT_REGISTERS_21_12_port);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => N674, CK => CLK, Q => 
                           n_1755, QN => n1396_port);
   NEXT_REGISTERS_reg_21_11_inst : DLH_X1 port map( G => n12076, D => N2896, Q 
                           => NEXT_REGISTERS_21_11_port);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => N673, CK => CLK, Q => 
                           n_1756, QN => n1397_port);
   NEXT_REGISTERS_reg_21_10_inst : DLH_X1 port map( G => n12076, D => N2895, Q 
                           => NEXT_REGISTERS_21_10_port);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => N672, CK => CLK, Q => 
                           n_1757, QN => n1398_port);
   NEXT_REGISTERS_reg_21_9_inst : DLH_X1 port map( G => n12076, D => N2894, Q 
                           => NEXT_REGISTERS_21_9_port);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => N671, CK => CLK, Q => n_1758
                           , QN => n1399_port);
   NEXT_REGISTERS_reg_21_8_inst : DLH_X1 port map( G => n12077, D => N2893, Q 
                           => NEXT_REGISTERS_21_8_port);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => N670, CK => CLK, Q => n_1759
                           , QN => n1400_port);
   NEXT_REGISTERS_reg_21_7_inst : DLH_X1 port map( G => n12077, D => N2892, Q 
                           => NEXT_REGISTERS_21_7_port);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => N669, CK => CLK, Q => n_1760
                           , QN => n1401_port);
   NEXT_REGISTERS_reg_21_6_inst : DLH_X1 port map( G => n12077, D => N2891, Q 
                           => NEXT_REGISTERS_21_6_port);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => N668, CK => CLK, Q => n_1761
                           , QN => n1402_port);
   NEXT_REGISTERS_reg_21_5_inst : DLH_X1 port map( G => n12077, D => N2890, Q 
                           => NEXT_REGISTERS_21_5_port);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => N667, CK => CLK, Q => n_1762
                           , QN => n1403_port);
   NEXT_REGISTERS_reg_21_4_inst : DLH_X1 port map( G => n12077, D => N2889, Q 
                           => NEXT_REGISTERS_21_4_port);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => N666, CK => CLK, Q => n_1763
                           , QN => n1404_port);
   NEXT_REGISTERS_reg_21_3_inst : DLH_X1 port map( G => n12077, D => N2888, Q 
                           => NEXT_REGISTERS_21_3_port);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => N665, CK => CLK, Q => n_1764
                           , QN => n1405_port);
   NEXT_REGISTERS_reg_21_2_inst : DLH_X1 port map( G => n12077, D => N2887, Q 
                           => NEXT_REGISTERS_21_2_port);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => N664, CK => CLK, Q => n_1765
                           , QN => n1406_port);
   NEXT_REGISTERS_reg_21_1_inst : DLH_X1 port map( G => n12077, D => N2886, Q 
                           => NEXT_REGISTERS_21_1_port);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => N663, CK => CLK, Q => n_1766
                           , QN => n1407_port);
   NEXT_REGISTERS_reg_21_0_inst : DLH_X1 port map( G => n12077, D => N2885, Q 
                           => NEXT_REGISTERS_21_0_port);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => N662, CK => CLK, Q => n_1767
                           , QN => n1408_port);
   NEXT_REGISTERS_reg_22_63_inst : DLH_X1 port map( G => n12081, D => N2883, Q 
                           => NEXT_REGISTERS_22_63_port);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => N661, CK => CLK, Q => 
                           n_1768, QN => n1409_port);
   NEXT_REGISTERS_reg_22_62_inst : DLH_X1 port map( G => n12081, D => N2882, Q 
                           => NEXT_REGISTERS_22_62_port);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => N660, CK => CLK, Q => 
                           n_1769, QN => n1410_port);
   NEXT_REGISTERS_reg_22_61_inst : DLH_X1 port map( G => n12081, D => N2881, Q 
                           => NEXT_REGISTERS_22_61_port);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => N659, CK => CLK, Q => 
                           n_1770, QN => n1411_port);
   NEXT_REGISTERS_reg_22_60_inst : DLH_X1 port map( G => n12081, D => N2880, Q 
                           => NEXT_REGISTERS_22_60_port);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => N658, CK => CLK, Q => 
                           n_1771, QN => n1412_port);
   NEXT_REGISTERS_reg_22_59_inst : DLH_X1 port map( G => n12081, D => N2879, Q 
                           => NEXT_REGISTERS_22_59_port);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => N657, CK => CLK, Q => 
                           n_1772, QN => n1413_port);
   NEXT_REGISTERS_reg_22_58_inst : DLH_X1 port map( G => n12081, D => N2878, Q 
                           => NEXT_REGISTERS_22_58_port);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => N656, CK => CLK, Q => 
                           n_1773, QN => n1414_port);
   NEXT_REGISTERS_reg_22_57_inst : DLH_X1 port map( G => n12081, D => N2877, Q 
                           => NEXT_REGISTERS_22_57_port);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => N655, CK => CLK, Q => 
                           n_1774, QN => n1415_port);
   NEXT_REGISTERS_reg_22_56_inst : DLH_X1 port map( G => n12081, D => N2876, Q 
                           => NEXT_REGISTERS_22_56_port);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => N654, CK => CLK, Q => 
                           n_1775, QN => n1416_port);
   NEXT_REGISTERS_reg_22_55_inst : DLH_X1 port map( G => n12081, D => N2875, Q 
                           => NEXT_REGISTERS_22_55_port);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => N653, CK => CLK, Q => 
                           n_1776, QN => n1417_port);
   NEXT_REGISTERS_reg_22_54_inst : DLH_X1 port map( G => n12081, D => N2874, Q 
                           => NEXT_REGISTERS_22_54_port);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => N652, CK => CLK, Q => 
                           n_1777, QN => n1418_port);
   NEXT_REGISTERS_reg_22_53_inst : DLH_X1 port map( G => n12081, D => N2873, Q 
                           => NEXT_REGISTERS_22_53_port);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => N651, CK => CLK, Q => 
                           n_1778, QN => n1419_port);
   NEXT_REGISTERS_reg_22_52_inst : DLH_X1 port map( G => n12082, D => N2872, Q 
                           => NEXT_REGISTERS_22_52_port);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => N650, CK => CLK, Q => 
                           n_1779, QN => n1420_port);
   NEXT_REGISTERS_reg_22_51_inst : DLH_X1 port map( G => n12082, D => N2871, Q 
                           => NEXT_REGISTERS_22_51_port);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => N649, CK => CLK, Q => 
                           n_1780, QN => n1421_port);
   NEXT_REGISTERS_reg_22_50_inst : DLH_X1 port map( G => n12082, D => N2870, Q 
                           => NEXT_REGISTERS_22_50_port);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => N648, CK => CLK, Q => 
                           n_1781, QN => n1422_port);
   NEXT_REGISTERS_reg_22_49_inst : DLH_X1 port map( G => n12082, D => N2869, Q 
                           => NEXT_REGISTERS_22_49_port);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => N647, CK => CLK, Q => 
                           n_1782, QN => n1423_port);
   NEXT_REGISTERS_reg_22_48_inst : DLH_X1 port map( G => n12082, D => N2868, Q 
                           => NEXT_REGISTERS_22_48_port);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => N646, CK => CLK, Q => 
                           n_1783, QN => n1424_port);
   NEXT_REGISTERS_reg_22_47_inst : DLH_X1 port map( G => n12082, D => N2867, Q 
                           => NEXT_REGISTERS_22_47_port);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => N645, CK => CLK, Q => 
                           n_1784, QN => n1425_port);
   NEXT_REGISTERS_reg_22_46_inst : DLH_X1 port map( G => n12082, D => N2866, Q 
                           => NEXT_REGISTERS_22_46_port);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => N644, CK => CLK, Q => 
                           n_1785, QN => n1426_port);
   NEXT_REGISTERS_reg_22_45_inst : DLH_X1 port map( G => n12082, D => N2865, Q 
                           => NEXT_REGISTERS_22_45_port);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => N643, CK => CLK, Q => 
                           n_1786, QN => n1427_port);
   NEXT_REGISTERS_reg_22_44_inst : DLH_X1 port map( G => n12082, D => N2864, Q 
                           => NEXT_REGISTERS_22_44_port);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => N642, CK => CLK, Q => 
                           n_1787, QN => n1428_port);
   NEXT_REGISTERS_reg_22_43_inst : DLH_X1 port map( G => n12082, D => N2863, Q 
                           => NEXT_REGISTERS_22_43_port);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => N641, CK => CLK, Q => 
                           n_1788, QN => n1429_port);
   NEXT_REGISTERS_reg_22_42_inst : DLH_X1 port map( G => n12082, D => N2862, Q 
                           => NEXT_REGISTERS_22_42_port);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => N640, CK => CLK, Q => 
                           n_1789, QN => n1430_port);
   NEXT_REGISTERS_reg_22_41_inst : DLH_X1 port map( G => n12083, D => N2861, Q 
                           => NEXT_REGISTERS_22_41_port);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => N639, CK => CLK, Q => 
                           n_1790, QN => n1431_port);
   NEXT_REGISTERS_reg_22_40_inst : DLH_X1 port map( G => n12083, D => N2860, Q 
                           => NEXT_REGISTERS_22_40_port);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => N638, CK => CLK, Q => 
                           n_1791, QN => n1432_port);
   NEXT_REGISTERS_reg_22_39_inst : DLH_X1 port map( G => n12083, D => N2859, Q 
                           => NEXT_REGISTERS_22_39_port);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => N637, CK => CLK, Q => 
                           n_1792, QN => n1433_port);
   NEXT_REGISTERS_reg_22_38_inst : DLH_X1 port map( G => n12083, D => N2858, Q 
                           => NEXT_REGISTERS_22_38_port);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => N636, CK => CLK, Q => 
                           n_1793, QN => n1434_port);
   NEXT_REGISTERS_reg_22_37_inst : DLH_X1 port map( G => n12083, D => N2857, Q 
                           => NEXT_REGISTERS_22_37_port);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => N635, CK => CLK, Q => 
                           n_1794, QN => n1435_port);
   NEXT_REGISTERS_reg_22_36_inst : DLH_X1 port map( G => n12083, D => N2856, Q 
                           => NEXT_REGISTERS_22_36_port);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => N634, CK => CLK, Q => 
                           n_1795, QN => n1436_port);
   NEXT_REGISTERS_reg_22_35_inst : DLH_X1 port map( G => n12083, D => N2855, Q 
                           => NEXT_REGISTERS_22_35_port);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => N633, CK => CLK, Q => 
                           n_1796, QN => n1437_port);
   NEXT_REGISTERS_reg_22_34_inst : DLH_X1 port map( G => n12083, D => N2854, Q 
                           => NEXT_REGISTERS_22_34_port);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => N632, CK => CLK, Q => 
                           n_1797, QN => n1438_port);
   NEXT_REGISTERS_reg_22_33_inst : DLH_X1 port map( G => n12083, D => N2853, Q 
                           => NEXT_REGISTERS_22_33_port);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => N631, CK => CLK, Q => 
                           n_1798, QN => n1439_port);
   NEXT_REGISTERS_reg_22_32_inst : DLH_X1 port map( G => n12083, D => N2852, Q 
                           => NEXT_REGISTERS_22_32_port);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => N630, CK => CLK, Q => 
                           n_1799, QN => n1440_port);
   NEXT_REGISTERS_reg_22_31_inst : DLH_X1 port map( G => n12083, D => N2851, Q 
                           => NEXT_REGISTERS_22_31_port);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => N629, CK => CLK, Q => 
                           n_1800, QN => n1441_port);
   NEXT_REGISTERS_reg_22_30_inst : DLH_X1 port map( G => n12084, D => N2850, Q 
                           => NEXT_REGISTERS_22_30_port);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => N628, CK => CLK, Q => 
                           n_1801, QN => n1442_port);
   NEXT_REGISTERS_reg_22_29_inst : DLH_X1 port map( G => n12084, D => N2849, Q 
                           => NEXT_REGISTERS_22_29_port);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => N627, CK => CLK, Q => 
                           n_1802, QN => n1443_port);
   NEXT_REGISTERS_reg_22_28_inst : DLH_X1 port map( G => n12084, D => N2848, Q 
                           => NEXT_REGISTERS_22_28_port);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => N626, CK => CLK, Q => 
                           n_1803, QN => n1444_port);
   NEXT_REGISTERS_reg_22_27_inst : DLH_X1 port map( G => n12084, D => N2847, Q 
                           => NEXT_REGISTERS_22_27_port);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => N625, CK => CLK, Q => 
                           n_1804, QN => n1445_port);
   NEXT_REGISTERS_reg_22_26_inst : DLH_X1 port map( G => n12084, D => N2846, Q 
                           => NEXT_REGISTERS_22_26_port);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => N624, CK => CLK, Q => 
                           n_1805, QN => n1446_port);
   NEXT_REGISTERS_reg_22_25_inst : DLH_X1 port map( G => n12084, D => N2845, Q 
                           => NEXT_REGISTERS_22_25_port);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => N623, CK => CLK, Q => 
                           n_1806, QN => n1447_port);
   NEXT_REGISTERS_reg_22_24_inst : DLH_X1 port map( G => n12084, D => N2844, Q 
                           => NEXT_REGISTERS_22_24_port);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => N622, CK => CLK, Q => 
                           n_1807, QN => n1448_port);
   NEXT_REGISTERS_reg_22_23_inst : DLH_X1 port map( G => n12084, D => N2843, Q 
                           => NEXT_REGISTERS_22_23_port);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => N621, CK => CLK, Q => 
                           n_1808, QN => n1449_port);
   NEXT_REGISTERS_reg_22_22_inst : DLH_X1 port map( G => n12084, D => N2842, Q 
                           => NEXT_REGISTERS_22_22_port);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => N620, CK => CLK, Q => 
                           n_1809, QN => n1450_port);
   NEXT_REGISTERS_reg_22_21_inst : DLH_X1 port map( G => n12084, D => N2841, Q 
                           => NEXT_REGISTERS_22_21_port);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => N619, CK => CLK, Q => 
                           n_1810, QN => n1451_port);
   NEXT_REGISTERS_reg_22_20_inst : DLH_X1 port map( G => n12084, D => N2840, Q 
                           => NEXT_REGISTERS_22_20_port);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => N618, CK => CLK, Q => 
                           n_1811, QN => n1452_port);
   NEXT_REGISTERS_reg_22_19_inst : DLH_X1 port map( G => n12085, D => N2839, Q 
                           => NEXT_REGISTERS_22_19_port);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => N617, CK => CLK, Q => 
                           n_1812, QN => n1453_port);
   NEXT_REGISTERS_reg_22_18_inst : DLH_X1 port map( G => n12085, D => N2838, Q 
                           => NEXT_REGISTERS_22_18_port);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => N616, CK => CLK, Q => 
                           n_1813, QN => n1454_port);
   NEXT_REGISTERS_reg_22_17_inst : DLH_X1 port map( G => n12085, D => N2837, Q 
                           => NEXT_REGISTERS_22_17_port);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => N615, CK => CLK, Q => 
                           n_1814, QN => n1455_port);
   NEXT_REGISTERS_reg_22_16_inst : DLH_X1 port map( G => n12085, D => N2836, Q 
                           => NEXT_REGISTERS_22_16_port);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => N614, CK => CLK, Q => 
                           n_1815, QN => n1456_port);
   NEXT_REGISTERS_reg_22_15_inst : DLH_X1 port map( G => n12085, D => N2835, Q 
                           => NEXT_REGISTERS_22_15_port);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => N613, CK => CLK, Q => 
                           n_1816, QN => n1457_port);
   NEXT_REGISTERS_reg_22_14_inst : DLH_X1 port map( G => n12085, D => N2834, Q 
                           => NEXT_REGISTERS_22_14_port);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => N612, CK => CLK, Q => 
                           n_1817, QN => n1458_port);
   NEXT_REGISTERS_reg_22_13_inst : DLH_X1 port map( G => n12085, D => N2833, Q 
                           => NEXT_REGISTERS_22_13_port);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => N611, CK => CLK, Q => 
                           n_1818, QN => n1459_port);
   NEXT_REGISTERS_reg_22_12_inst : DLH_X1 port map( G => n12085, D => N2832, Q 
                           => NEXT_REGISTERS_22_12_port);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => N610, CK => CLK, Q => 
                           n_1819, QN => n1460_port);
   NEXT_REGISTERS_reg_22_11_inst : DLH_X1 port map( G => n12085, D => N2831, Q 
                           => NEXT_REGISTERS_22_11_port);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => N609, CK => CLK, Q => 
                           n_1820, QN => n1461_port);
   NEXT_REGISTERS_reg_22_10_inst : DLH_X1 port map( G => n12085, D => N2830, Q 
                           => NEXT_REGISTERS_22_10_port);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => N608, CK => CLK, Q => 
                           n_1821, QN => n1462_port);
   NEXT_REGISTERS_reg_22_9_inst : DLH_X1 port map( G => n12085, D => N2829, Q 
                           => NEXT_REGISTERS_22_9_port);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => N607, CK => CLK, Q => n_1822
                           , QN => n1463_port);
   NEXT_REGISTERS_reg_22_8_inst : DLH_X1 port map( G => n12086, D => N2828, Q 
                           => NEXT_REGISTERS_22_8_port);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => N606, CK => CLK, Q => n_1823
                           , QN => n1464_port);
   NEXT_REGISTERS_reg_22_7_inst : DLH_X1 port map( G => n12086, D => N2827, Q 
                           => NEXT_REGISTERS_22_7_port);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => N605, CK => CLK, Q => n_1824
                           , QN => n1465_port);
   NEXT_REGISTERS_reg_22_6_inst : DLH_X1 port map( G => n12086, D => N2826, Q 
                           => NEXT_REGISTERS_22_6_port);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => N604, CK => CLK, Q => n_1825
                           , QN => n1466_port);
   NEXT_REGISTERS_reg_22_5_inst : DLH_X1 port map( G => n12086, D => N2825, Q 
                           => NEXT_REGISTERS_22_5_port);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => N603, CK => CLK, Q => n_1826
                           , QN => n1467_port);
   NEXT_REGISTERS_reg_22_4_inst : DLH_X1 port map( G => n12086, D => N2824, Q 
                           => NEXT_REGISTERS_22_4_port);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => N602, CK => CLK, Q => n_1827
                           , QN => n1468_port);
   NEXT_REGISTERS_reg_22_3_inst : DLH_X1 port map( G => n12086, D => N2823, Q 
                           => NEXT_REGISTERS_22_3_port);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => N601, CK => CLK, Q => n_1828
                           , QN => n1469_port);
   NEXT_REGISTERS_reg_22_2_inst : DLH_X1 port map( G => n12086, D => N2822, Q 
                           => NEXT_REGISTERS_22_2_port);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => N600, CK => CLK, Q => n_1829
                           , QN => n1470_port);
   NEXT_REGISTERS_reg_22_1_inst : DLH_X1 port map( G => n12086, D => N2821, Q 
                           => NEXT_REGISTERS_22_1_port);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => N599, CK => CLK, Q => n_1830
                           , QN => n1471_port);
   NEXT_REGISTERS_reg_22_0_inst : DLH_X1 port map( G => n12086, D => N2820, Q 
                           => NEXT_REGISTERS_22_0_port);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => N598, CK => CLK, Q => n_1831
                           , QN => n1472_port);
   NEXT_REGISTERS_reg_23_63_inst : DLH_X1 port map( G => n12090, D => N2818, Q 
                           => NEXT_REGISTERS_23_63_port);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => N597, CK => CLK, Q => 
                           n10285, QN => n1473_port);
   NEXT_REGISTERS_reg_23_62_inst : DLH_X1 port map( G => n12090, D => N2817, Q 
                           => NEXT_REGISTERS_23_62_port);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => N596, CK => CLK, Q => 
                           n10283, QN => n1474_port);
   NEXT_REGISTERS_reg_23_61_inst : DLH_X1 port map( G => n12090, D => N2816, Q 
                           => NEXT_REGISTERS_23_61_port);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => N595, CK => CLK, Q => 
                           n10281, QN => n1475_port);
   NEXT_REGISTERS_reg_23_60_inst : DLH_X1 port map( G => n12090, D => N2815, Q 
                           => NEXT_REGISTERS_23_60_port);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => N594, CK => CLK, Q => 
                           n10279, QN => n1476_port);
   NEXT_REGISTERS_reg_23_59_inst : DLH_X1 port map( G => n12090, D => N2814, Q 
                           => NEXT_REGISTERS_23_59_port);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => N593, CK => CLK, Q => 
                           n10277, QN => n1477_port);
   NEXT_REGISTERS_reg_23_58_inst : DLH_X1 port map( G => n12090, D => N2813, Q 
                           => NEXT_REGISTERS_23_58_port);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => N592, CK => CLK, Q => 
                           n10275, QN => n1478_port);
   NEXT_REGISTERS_reg_23_57_inst : DLH_X1 port map( G => n12090, D => N2812, Q 
                           => NEXT_REGISTERS_23_57_port);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => N591, CK => CLK, Q => 
                           n10273, QN => n1479_port);
   NEXT_REGISTERS_reg_23_56_inst : DLH_X1 port map( G => n12090, D => N2811, Q 
                           => NEXT_REGISTERS_23_56_port);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => N590, CK => CLK, Q => 
                           n10271, QN => n1480_port);
   NEXT_REGISTERS_reg_23_55_inst : DLH_X1 port map( G => n12090, D => N2810, Q 
                           => NEXT_REGISTERS_23_55_port);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => N589, CK => CLK, Q => 
                           n10269, QN => n1481_port);
   NEXT_REGISTERS_reg_23_54_inst : DLH_X1 port map( G => n12090, D => N2809, Q 
                           => NEXT_REGISTERS_23_54_port);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => N588, CK => CLK, Q => 
                           n10267, QN => n1482_port);
   NEXT_REGISTERS_reg_23_53_inst : DLH_X1 port map( G => n12090, D => N2808, Q 
                           => NEXT_REGISTERS_23_53_port);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => N587, CK => CLK, Q => 
                           n10265, QN => n1483_port);
   NEXT_REGISTERS_reg_23_52_inst : DLH_X1 port map( G => n12091, D => N2807, Q 
                           => NEXT_REGISTERS_23_52_port);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => N586, CK => CLK, Q => 
                           n10263, QN => n1484_port);
   NEXT_REGISTERS_reg_23_51_inst : DLH_X1 port map( G => n12091, D => N2806, Q 
                           => NEXT_REGISTERS_23_51_port);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => N585, CK => CLK, Q => 
                           n10261, QN => n1485_port);
   NEXT_REGISTERS_reg_23_50_inst : DLH_X1 port map( G => n12091, D => N2805, Q 
                           => NEXT_REGISTERS_23_50_port);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => N584, CK => CLK, Q => 
                           n10259, QN => n1486_port);
   NEXT_REGISTERS_reg_23_49_inst : DLH_X1 port map( G => n12091, D => N2804, Q 
                           => NEXT_REGISTERS_23_49_port);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => N583, CK => CLK, Q => 
                           n10257, QN => n1487_port);
   NEXT_REGISTERS_reg_23_48_inst : DLH_X1 port map( G => n12091, D => N2803, Q 
                           => NEXT_REGISTERS_23_48_port);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => N582, CK => CLK, Q => 
                           n10255, QN => n1488_port);
   NEXT_REGISTERS_reg_23_47_inst : DLH_X1 port map( G => n12091, D => N2802, Q 
                           => NEXT_REGISTERS_23_47_port);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => N581, CK => CLK, Q => 
                           n10253, QN => n1489_port);
   NEXT_REGISTERS_reg_23_46_inst : DLH_X1 port map( G => n12091, D => N2801, Q 
                           => NEXT_REGISTERS_23_46_port);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => N580, CK => CLK, Q => 
                           n10251, QN => n1490_port);
   NEXT_REGISTERS_reg_23_45_inst : DLH_X1 port map( G => n12091, D => N2800, Q 
                           => NEXT_REGISTERS_23_45_port);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => N579, CK => CLK, Q => 
                           n10249, QN => n1491_port);
   NEXT_REGISTERS_reg_23_44_inst : DLH_X1 port map( G => n12091, D => N2799, Q 
                           => NEXT_REGISTERS_23_44_port);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => N578, CK => CLK, Q => 
                           n10247, QN => n1492_port);
   NEXT_REGISTERS_reg_23_43_inst : DLH_X1 port map( G => n12091, D => N2798, Q 
                           => NEXT_REGISTERS_23_43_port);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => N577, CK => CLK, Q => 
                           n10245, QN => n1493_port);
   NEXT_REGISTERS_reg_23_42_inst : DLH_X1 port map( G => n12091, D => N2797, Q 
                           => NEXT_REGISTERS_23_42_port);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => N576, CK => CLK, Q => 
                           n10243, QN => n1494_port);
   NEXT_REGISTERS_reg_23_41_inst : DLH_X1 port map( G => n12092, D => N2796, Q 
                           => NEXT_REGISTERS_23_41_port);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => N575, CK => CLK, Q => 
                           n10241, QN => n1495_port);
   NEXT_REGISTERS_reg_23_40_inst : DLH_X1 port map( G => n12092, D => N2795, Q 
                           => NEXT_REGISTERS_23_40_port);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => N574, CK => CLK, Q => 
                           n10239, QN => n1496_port);
   NEXT_REGISTERS_reg_23_39_inst : DLH_X1 port map( G => n12092, D => N2794, Q 
                           => NEXT_REGISTERS_23_39_port);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => N573, CK => CLK, Q => 
                           n10237, QN => n1497_port);
   NEXT_REGISTERS_reg_23_38_inst : DLH_X1 port map( G => n12092, D => N2793, Q 
                           => NEXT_REGISTERS_23_38_port);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => N572, CK => CLK, Q => 
                           n10235, QN => n1498_port);
   NEXT_REGISTERS_reg_23_37_inst : DLH_X1 port map( G => n12092, D => N2792, Q 
                           => NEXT_REGISTERS_23_37_port);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => N571, CK => CLK, Q => 
                           n10233, QN => n1499_port);
   NEXT_REGISTERS_reg_23_36_inst : DLH_X1 port map( G => n12092, D => N2791, Q 
                           => NEXT_REGISTERS_23_36_port);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => N570, CK => CLK, Q => 
                           n10231, QN => n1500_port);
   NEXT_REGISTERS_reg_23_35_inst : DLH_X1 port map( G => n12092, D => N2790, Q 
                           => NEXT_REGISTERS_23_35_port);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => N569, CK => CLK, Q => 
                           n10229, QN => n1501_port);
   NEXT_REGISTERS_reg_23_34_inst : DLH_X1 port map( G => n12092, D => N2789, Q 
                           => NEXT_REGISTERS_23_34_port);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => N568, CK => CLK, Q => 
                           n10227, QN => n1502_port);
   NEXT_REGISTERS_reg_23_33_inst : DLH_X1 port map( G => n12092, D => N2788, Q 
                           => NEXT_REGISTERS_23_33_port);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => N567, CK => CLK, Q => 
                           n10225, QN => n1503_port);
   NEXT_REGISTERS_reg_23_32_inst : DLH_X1 port map( G => n12092, D => N2787, Q 
                           => NEXT_REGISTERS_23_32_port);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => N566, CK => CLK, Q => 
                           n10223, QN => n1504_port);
   NEXT_REGISTERS_reg_23_31_inst : DLH_X1 port map( G => n12092, D => N2786, Q 
                           => NEXT_REGISTERS_23_31_port);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => N565, CK => CLK, Q => 
                           n10221, QN => n1505_port);
   NEXT_REGISTERS_reg_23_30_inst : DLH_X1 port map( G => n12093, D => N2785, Q 
                           => NEXT_REGISTERS_23_30_port);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => N564, CK => CLK, Q => 
                           n10219, QN => n1506_port);
   NEXT_REGISTERS_reg_23_29_inst : DLH_X1 port map( G => n12093, D => N2784, Q 
                           => NEXT_REGISTERS_23_29_port);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => N563, CK => CLK, Q => 
                           n10217, QN => n1507_port);
   NEXT_REGISTERS_reg_23_28_inst : DLH_X1 port map( G => n12093, D => N2783, Q 
                           => NEXT_REGISTERS_23_28_port);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => N562, CK => CLK, Q => 
                           n10215, QN => n1508_port);
   NEXT_REGISTERS_reg_23_27_inst : DLH_X1 port map( G => n12093, D => N2782, Q 
                           => NEXT_REGISTERS_23_27_port);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => N561, CK => CLK, Q => 
                           n10213, QN => n1509_port);
   NEXT_REGISTERS_reg_23_26_inst : DLH_X1 port map( G => n12093, D => N2781, Q 
                           => NEXT_REGISTERS_23_26_port);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => N560, CK => CLK, Q => 
                           n10211, QN => n1510_port);
   NEXT_REGISTERS_reg_23_25_inst : DLH_X1 port map( G => n12093, D => N2780, Q 
                           => NEXT_REGISTERS_23_25_port);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => N559, CK => CLK, Q => 
                           n10209, QN => n1511_port);
   NEXT_REGISTERS_reg_23_24_inst : DLH_X1 port map( G => n12093, D => N2779, Q 
                           => NEXT_REGISTERS_23_24_port);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => N558, CK => CLK, Q => 
                           n10207, QN => n1512_port);
   NEXT_REGISTERS_reg_23_23_inst : DLH_X1 port map( G => n12093, D => N2778, Q 
                           => NEXT_REGISTERS_23_23_port);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => N557, CK => CLK, Q => 
                           n10205, QN => n1513_port);
   NEXT_REGISTERS_reg_23_22_inst : DLH_X1 port map( G => n12093, D => N2777, Q 
                           => NEXT_REGISTERS_23_22_port);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => N556, CK => CLK, Q => 
                           n10203, QN => n1514_port);
   NEXT_REGISTERS_reg_23_21_inst : DLH_X1 port map( G => n12093, D => N2776, Q 
                           => NEXT_REGISTERS_23_21_port);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => N555, CK => CLK, Q => 
                           n10201, QN => n1515_port);
   NEXT_REGISTERS_reg_23_20_inst : DLH_X1 port map( G => n12093, D => N2775, Q 
                           => NEXT_REGISTERS_23_20_port);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => N554, CK => CLK, Q => 
                           n10199, QN => n1516_port);
   NEXT_REGISTERS_reg_23_19_inst : DLH_X1 port map( G => n12094, D => N2774, Q 
                           => NEXT_REGISTERS_23_19_port);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => N553, CK => CLK, Q => 
                           n10197, QN => n1517_port);
   NEXT_REGISTERS_reg_23_18_inst : DLH_X1 port map( G => n12094, D => N2773, Q 
                           => NEXT_REGISTERS_23_18_port);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => N552, CK => CLK, Q => 
                           n10195, QN => n1518_port);
   NEXT_REGISTERS_reg_23_17_inst : DLH_X1 port map( G => n12094, D => N2772, Q 
                           => NEXT_REGISTERS_23_17_port);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => N551, CK => CLK, Q => 
                           n10193, QN => n1519_port);
   NEXT_REGISTERS_reg_23_16_inst : DLH_X1 port map( G => n12094, D => N2771, Q 
                           => NEXT_REGISTERS_23_16_port);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => N550, CK => CLK, Q => 
                           n10191, QN => n1520_port);
   NEXT_REGISTERS_reg_23_15_inst : DLH_X1 port map( G => n12094, D => N2770, Q 
                           => NEXT_REGISTERS_23_15_port);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => N549, CK => CLK, Q => 
                           n10189, QN => n1521_port);
   NEXT_REGISTERS_reg_23_14_inst : DLH_X1 port map( G => n12094, D => N2769, Q 
                           => NEXT_REGISTERS_23_14_port);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => N548, CK => CLK, Q => 
                           n10187, QN => n1522_port);
   NEXT_REGISTERS_reg_23_13_inst : DLH_X1 port map( G => n12094, D => N2768, Q 
                           => NEXT_REGISTERS_23_13_port);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => N547, CK => CLK, Q => 
                           n10185, QN => n1523_port);
   NEXT_REGISTERS_reg_23_12_inst : DLH_X1 port map( G => n12094, D => N2767, Q 
                           => NEXT_REGISTERS_23_12_port);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => N546, CK => CLK, Q => 
                           n10183, QN => n1524_port);
   NEXT_REGISTERS_reg_23_11_inst : DLH_X1 port map( G => n12094, D => N2766, Q 
                           => NEXT_REGISTERS_23_11_port);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => N545, CK => CLK, Q => 
                           n10181, QN => n1525_port);
   NEXT_REGISTERS_reg_23_10_inst : DLH_X1 port map( G => n12094, D => N2765, Q 
                           => NEXT_REGISTERS_23_10_port);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => N544, CK => CLK, Q => 
                           n10179, QN => n1526_port);
   NEXT_REGISTERS_reg_23_9_inst : DLH_X1 port map( G => n12094, D => N2764, Q 
                           => NEXT_REGISTERS_23_9_port);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => N543, CK => CLK, Q => n10177
                           , QN => n1527_port);
   NEXT_REGISTERS_reg_23_8_inst : DLH_X1 port map( G => n12095, D => N2763, Q 
                           => NEXT_REGISTERS_23_8_port);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => N542, CK => CLK, Q => n10175
                           , QN => n1528_port);
   NEXT_REGISTERS_reg_23_7_inst : DLH_X1 port map( G => n12095, D => N2762, Q 
                           => NEXT_REGISTERS_23_7_port);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => N541, CK => CLK, Q => n10173
                           , QN => n1529_port);
   NEXT_REGISTERS_reg_23_6_inst : DLH_X1 port map( G => n12095, D => N2761, Q 
                           => NEXT_REGISTERS_23_6_port);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => N540, CK => CLK, Q => n10171
                           , QN => n1530_port);
   NEXT_REGISTERS_reg_23_5_inst : DLH_X1 port map( G => n12095, D => N2760, Q 
                           => NEXT_REGISTERS_23_5_port);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => N539, CK => CLK, Q => n10169
                           , QN => n1531_port);
   NEXT_REGISTERS_reg_23_4_inst : DLH_X1 port map( G => n12095, D => N2759, Q 
                           => NEXT_REGISTERS_23_4_port);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => N538, CK => CLK, Q => n10167
                           , QN => n1532_port);
   NEXT_REGISTERS_reg_23_3_inst : DLH_X1 port map( G => n12095, D => N2758, Q 
                           => NEXT_REGISTERS_23_3_port);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => N537, CK => CLK, Q => n10165
                           , QN => n1533_port);
   NEXT_REGISTERS_reg_23_2_inst : DLH_X1 port map( G => n12095, D => N2757, Q 
                           => NEXT_REGISTERS_23_2_port);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => N536, CK => CLK, Q => n10163
                           , QN => n1534_port);
   NEXT_REGISTERS_reg_23_1_inst : DLH_X1 port map( G => n12095, D => N2756, Q 
                           => NEXT_REGISTERS_23_1_port);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => N535, CK => CLK, Q => n10161
                           , QN => n1535_port);
   NEXT_REGISTERS_reg_23_0_inst : DLH_X1 port map( G => n12095, D => N2755, Q 
                           => NEXT_REGISTERS_23_0_port);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => N534, CK => CLK, Q => n10159
                           , QN => n1536_port);
   NEXT_REGISTERS_reg_24_63_inst : DLH_X1 port map( G => n12099, D => N2753, Q 
                           => NEXT_REGISTERS_24_63_port);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => N533, CK => CLK, Q => n9837
                           , QN => n1537_port);
   NEXT_REGISTERS_reg_24_62_inst : DLH_X1 port map( G => n12099, D => N2752, Q 
                           => NEXT_REGISTERS_24_62_port);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => N532, CK => CLK, Q => n9835
                           , QN => n1538_port);
   NEXT_REGISTERS_reg_24_61_inst : DLH_X1 port map( G => n12099, D => N2751, Q 
                           => NEXT_REGISTERS_24_61_port);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => N531, CK => CLK, Q => n9833
                           , QN => n1539_port);
   NEXT_REGISTERS_reg_24_60_inst : DLH_X1 port map( G => n12099, D => N2750, Q 
                           => NEXT_REGISTERS_24_60_port);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => N530, CK => CLK, Q => n9831
                           , QN => n1540_port);
   NEXT_REGISTERS_reg_24_59_inst : DLH_X1 port map( G => n12099, D => N2749, Q 
                           => NEXT_REGISTERS_24_59_port);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => N529, CK => CLK, Q => n9829
                           , QN => n1541_port);
   NEXT_REGISTERS_reg_24_58_inst : DLH_X1 port map( G => n12099, D => N2748, Q 
                           => NEXT_REGISTERS_24_58_port);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => N528, CK => CLK, Q => n9827
                           , QN => n1542_port);
   NEXT_REGISTERS_reg_24_57_inst : DLH_X1 port map( G => n12099, D => N2747, Q 
                           => NEXT_REGISTERS_24_57_port);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => N527, CK => CLK, Q => n9825
                           , QN => n1543_port);
   NEXT_REGISTERS_reg_24_56_inst : DLH_X1 port map( G => n12099, D => N2746, Q 
                           => NEXT_REGISTERS_24_56_port);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => N526, CK => CLK, Q => n9823
                           , QN => n1544_port);
   NEXT_REGISTERS_reg_24_55_inst : DLH_X1 port map( G => n12099, D => N2745, Q 
                           => NEXT_REGISTERS_24_55_port);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => N525, CK => CLK, Q => n9821
                           , QN => n1545_port);
   NEXT_REGISTERS_reg_24_54_inst : DLH_X1 port map( G => n12099, D => N2744, Q 
                           => NEXT_REGISTERS_24_54_port);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => N524, CK => CLK, Q => n9819
                           , QN => n1546_port);
   NEXT_REGISTERS_reg_24_53_inst : DLH_X1 port map( G => n12099, D => N2743, Q 
                           => NEXT_REGISTERS_24_53_port);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => N523, CK => CLK, Q => n9817
                           , QN => n1547_port);
   NEXT_REGISTERS_reg_24_52_inst : DLH_X1 port map( G => n12100, D => N2742, Q 
                           => NEXT_REGISTERS_24_52_port);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => N522, CK => CLK, Q => n9815
                           , QN => n1548_port);
   NEXT_REGISTERS_reg_24_51_inst : DLH_X1 port map( G => n12100, D => N2741, Q 
                           => NEXT_REGISTERS_24_51_port);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => N521, CK => CLK, Q => n9813
                           , QN => n1549_port);
   NEXT_REGISTERS_reg_24_50_inst : DLH_X1 port map( G => n12100, D => N2740, Q 
                           => NEXT_REGISTERS_24_50_port);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => N520, CK => CLK, Q => n9811
                           , QN => n1550_port);
   NEXT_REGISTERS_reg_24_49_inst : DLH_X1 port map( G => n12100, D => N2739, Q 
                           => NEXT_REGISTERS_24_49_port);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => N519, CK => CLK, Q => n9809
                           , QN => n1551_port);
   NEXT_REGISTERS_reg_24_48_inst : DLH_X1 port map( G => n12100, D => N2738, Q 
                           => NEXT_REGISTERS_24_48_port);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => N518, CK => CLK, Q => n9807
                           , QN => n1552_port);
   NEXT_REGISTERS_reg_24_47_inst : DLH_X1 port map( G => n12100, D => N2737, Q 
                           => NEXT_REGISTERS_24_47_port);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => N517, CK => CLK, Q => n9805
                           , QN => n1553_port);
   NEXT_REGISTERS_reg_24_46_inst : DLH_X1 port map( G => n12100, D => N2736, Q 
                           => NEXT_REGISTERS_24_46_port);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => N516, CK => CLK, Q => n9803
                           , QN => n1554_port);
   NEXT_REGISTERS_reg_24_45_inst : DLH_X1 port map( G => n12100, D => N2735, Q 
                           => NEXT_REGISTERS_24_45_port);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => N515, CK => CLK, Q => n9801
                           , QN => n1555_port);
   NEXT_REGISTERS_reg_24_44_inst : DLH_X1 port map( G => n12100, D => N2734, Q 
                           => NEXT_REGISTERS_24_44_port);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => N514, CK => CLK, Q => n9799
                           , QN => n1556_port);
   NEXT_REGISTERS_reg_24_43_inst : DLH_X1 port map( G => n12100, D => N2733, Q 
                           => NEXT_REGISTERS_24_43_port);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => N513, CK => CLK, Q => n9797
                           , QN => n1557_port);
   NEXT_REGISTERS_reg_24_42_inst : DLH_X1 port map( G => n12100, D => N2732, Q 
                           => NEXT_REGISTERS_24_42_port);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => N512, CK => CLK, Q => n9795
                           , QN => n1558_port);
   NEXT_REGISTERS_reg_24_41_inst : DLH_X1 port map( G => n12101, D => N2731, Q 
                           => NEXT_REGISTERS_24_41_port);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => N511, CK => CLK, Q => n9793
                           , QN => n1559_port);
   NEXT_REGISTERS_reg_24_40_inst : DLH_X1 port map( G => n12101, D => N2730, Q 
                           => NEXT_REGISTERS_24_40_port);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => N510, CK => CLK, Q => n9791
                           , QN => n1560_port);
   NEXT_REGISTERS_reg_24_39_inst : DLH_X1 port map( G => n12101, D => N2729, Q 
                           => NEXT_REGISTERS_24_39_port);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => N509, CK => CLK, Q => n9789
                           , QN => n1561_port);
   NEXT_REGISTERS_reg_24_38_inst : DLH_X1 port map( G => n12101, D => N2728, Q 
                           => NEXT_REGISTERS_24_38_port);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => N508, CK => CLK, Q => n9787
                           , QN => n1562_port);
   NEXT_REGISTERS_reg_24_37_inst : DLH_X1 port map( G => n12101, D => N2727, Q 
                           => NEXT_REGISTERS_24_37_port);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => N507, CK => CLK, Q => n9785
                           , QN => n1563_port);
   NEXT_REGISTERS_reg_24_36_inst : DLH_X1 port map( G => n12101, D => N2726, Q 
                           => NEXT_REGISTERS_24_36_port);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => N506, CK => CLK, Q => n9783
                           , QN => n1564_port);
   NEXT_REGISTERS_reg_24_35_inst : DLH_X1 port map( G => n12101, D => N2725, Q 
                           => NEXT_REGISTERS_24_35_port);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => N505, CK => CLK, Q => n9781
                           , QN => n1565_port);
   NEXT_REGISTERS_reg_24_34_inst : DLH_X1 port map( G => n12101, D => N2724, Q 
                           => NEXT_REGISTERS_24_34_port);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => N504, CK => CLK, Q => n9779
                           , QN => n1566_port);
   NEXT_REGISTERS_reg_24_33_inst : DLH_X1 port map( G => n12101, D => N2723, Q 
                           => NEXT_REGISTERS_24_33_port);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => N503, CK => CLK, Q => n9777
                           , QN => n1567_port);
   NEXT_REGISTERS_reg_24_32_inst : DLH_X1 port map( G => n12101, D => N2722, Q 
                           => NEXT_REGISTERS_24_32_port);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => N502, CK => CLK, Q => n9775
                           , QN => n1568_port);
   NEXT_REGISTERS_reg_24_31_inst : DLH_X1 port map( G => n12101, D => N2721, Q 
                           => NEXT_REGISTERS_24_31_port);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => N501, CK => CLK, Q => n9773
                           , QN => n1569_port);
   NEXT_REGISTERS_reg_24_30_inst : DLH_X1 port map( G => n12102, D => N2720, Q 
                           => NEXT_REGISTERS_24_30_port);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => N500, CK => CLK, Q => n9771
                           , QN => n1570_port);
   NEXT_REGISTERS_reg_24_29_inst : DLH_X1 port map( G => n12102, D => N2719, Q 
                           => NEXT_REGISTERS_24_29_port);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => N499, CK => CLK, Q => n9769
                           , QN => n1571_port);
   NEXT_REGISTERS_reg_24_28_inst : DLH_X1 port map( G => n12102, D => N2718, Q 
                           => NEXT_REGISTERS_24_28_port);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => N498, CK => CLK, Q => n9767
                           , QN => n1572_port);
   NEXT_REGISTERS_reg_24_27_inst : DLH_X1 port map( G => n12102, D => N2717, Q 
                           => NEXT_REGISTERS_24_27_port);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => N497, CK => CLK, Q => n9765
                           , QN => n1573_port);
   NEXT_REGISTERS_reg_24_26_inst : DLH_X1 port map( G => n12102, D => N2716, Q 
                           => NEXT_REGISTERS_24_26_port);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => N496, CK => CLK, Q => n9763
                           , QN => n1574_port);
   NEXT_REGISTERS_reg_24_25_inst : DLH_X1 port map( G => n12102, D => N2715, Q 
                           => NEXT_REGISTERS_24_25_port);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => N495, CK => CLK, Q => n9761
                           , QN => n1575_port);
   NEXT_REGISTERS_reg_24_24_inst : DLH_X1 port map( G => n12102, D => N2714, Q 
                           => NEXT_REGISTERS_24_24_port);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => N494, CK => CLK, Q => n9759
                           , QN => n1576_port);
   NEXT_REGISTERS_reg_24_23_inst : DLH_X1 port map( G => n12102, D => N2713, Q 
                           => NEXT_REGISTERS_24_23_port);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => N493, CK => CLK, Q => n9757
                           , QN => n1577_port);
   NEXT_REGISTERS_reg_24_22_inst : DLH_X1 port map( G => n12102, D => N2712, Q 
                           => NEXT_REGISTERS_24_22_port);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => N492, CK => CLK, Q => n9755
                           , QN => n1578_port);
   NEXT_REGISTERS_reg_24_21_inst : DLH_X1 port map( G => n12102, D => N2711, Q 
                           => NEXT_REGISTERS_24_21_port);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => N491, CK => CLK, Q => n9753
                           , QN => n1579_port);
   NEXT_REGISTERS_reg_24_20_inst : DLH_X1 port map( G => n12102, D => N2710, Q 
                           => NEXT_REGISTERS_24_20_port);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => N490, CK => CLK, Q => n9751
                           , QN => n1580_port);
   NEXT_REGISTERS_reg_24_19_inst : DLH_X1 port map( G => n12103, D => N2709, Q 
                           => NEXT_REGISTERS_24_19_port);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => N489, CK => CLK, Q => n9749
                           , QN => n1581_port);
   NEXT_REGISTERS_reg_24_18_inst : DLH_X1 port map( G => n12103, D => N2708, Q 
                           => NEXT_REGISTERS_24_18_port);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => N488, CK => CLK, Q => n9747
                           , QN => n1582_port);
   NEXT_REGISTERS_reg_24_17_inst : DLH_X1 port map( G => n12103, D => N2707, Q 
                           => NEXT_REGISTERS_24_17_port);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => N487, CK => CLK, Q => n9745
                           , QN => n1583_port);
   NEXT_REGISTERS_reg_24_16_inst : DLH_X1 port map( G => n12103, D => N2706, Q 
                           => NEXT_REGISTERS_24_16_port);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => N486, CK => CLK, Q => n9743
                           , QN => n1584_port);
   NEXT_REGISTERS_reg_24_15_inst : DLH_X1 port map( G => n12103, D => N2705, Q 
                           => NEXT_REGISTERS_24_15_port);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => N485, CK => CLK, Q => n9741
                           , QN => n1585_port);
   NEXT_REGISTERS_reg_24_14_inst : DLH_X1 port map( G => n12103, D => N2704, Q 
                           => NEXT_REGISTERS_24_14_port);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => N484, CK => CLK, Q => n9739
                           , QN => n1586_port);
   NEXT_REGISTERS_reg_24_13_inst : DLH_X1 port map( G => n12103, D => N2703, Q 
                           => NEXT_REGISTERS_24_13_port);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => N483, CK => CLK, Q => n9737
                           , QN => n1587_port);
   NEXT_REGISTERS_reg_24_12_inst : DLH_X1 port map( G => n12103, D => N2702, Q 
                           => NEXT_REGISTERS_24_12_port);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => N482, CK => CLK, Q => n9735
                           , QN => n1588_port);
   NEXT_REGISTERS_reg_24_11_inst : DLH_X1 port map( G => n12103, D => N2701, Q 
                           => NEXT_REGISTERS_24_11_port);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => N481, CK => CLK, Q => n9733
                           , QN => n1589_port);
   NEXT_REGISTERS_reg_24_10_inst : DLH_X1 port map( G => n12103, D => N2700, Q 
                           => NEXT_REGISTERS_24_10_port);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => N480, CK => CLK, Q => n9731
                           , QN => n1590_port);
   NEXT_REGISTERS_reg_24_9_inst : DLH_X1 port map( G => n12103, D => N2699, Q 
                           => NEXT_REGISTERS_24_9_port);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => N479, CK => CLK, Q => n9729,
                           QN => n1591_port);
   NEXT_REGISTERS_reg_24_8_inst : DLH_X1 port map( G => n12104, D => N2698, Q 
                           => NEXT_REGISTERS_24_8_port);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => N478, CK => CLK, Q => n9727,
                           QN => n1592_port);
   NEXT_REGISTERS_reg_24_7_inst : DLH_X1 port map( G => n12104, D => N2697, Q 
                           => NEXT_REGISTERS_24_7_port);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => N477, CK => CLK, Q => n9725,
                           QN => n1593_port);
   NEXT_REGISTERS_reg_24_6_inst : DLH_X1 port map( G => n12104, D => N2696, Q 
                           => NEXT_REGISTERS_24_6_port);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => N476, CK => CLK, Q => n9723,
                           QN => n1594_port);
   NEXT_REGISTERS_reg_24_5_inst : DLH_X1 port map( G => n12104, D => N2695, Q 
                           => NEXT_REGISTERS_24_5_port);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => N475, CK => CLK, Q => n9721,
                           QN => n1595_port);
   NEXT_REGISTERS_reg_24_4_inst : DLH_X1 port map( G => n12104, D => N2694, Q 
                           => NEXT_REGISTERS_24_4_port);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => N474, CK => CLK, Q => n9719,
                           QN => n1596_port);
   NEXT_REGISTERS_reg_24_3_inst : DLH_X1 port map( G => n12104, D => N2693, Q 
                           => NEXT_REGISTERS_24_3_port);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => N473, CK => CLK, Q => n9717,
                           QN => n1597_port);
   NEXT_REGISTERS_reg_24_2_inst : DLH_X1 port map( G => n12104, D => N2692, Q 
                           => NEXT_REGISTERS_24_2_port);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => N472, CK => CLK, Q => n9715,
                           QN => n1598_port);
   NEXT_REGISTERS_reg_24_1_inst : DLH_X1 port map( G => n12104, D => N2691, Q 
                           => NEXT_REGISTERS_24_1_port);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => N471, CK => CLK, Q => n9713,
                           QN => n1599_port);
   NEXT_REGISTERS_reg_24_0_inst : DLH_X1 port map( G => n12104, D => N2690, Q 
                           => NEXT_REGISTERS_24_0_port);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => N470, CK => CLK, Q => n9711,
                           QN => n1600_port);
   NEXT_REGISTERS_reg_25_63_inst : DLH_X1 port map( G => n12108, D => N2688, Q 
                           => NEXT_REGISTERS_25_63_port);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => N469, CK => CLK, Q => 
                           n10158, QN => n1601_port);
   NEXT_REGISTERS_reg_25_62_inst : DLH_X1 port map( G => n12108, D => N2687, Q 
                           => NEXT_REGISTERS_25_62_port);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => N468, CK => CLK, Q => 
                           n10157, QN => n1602_port);
   NEXT_REGISTERS_reg_25_61_inst : DLH_X1 port map( G => n12108, D => N2686, Q 
                           => NEXT_REGISTERS_25_61_port);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => N467, CK => CLK, Q => 
                           n10156, QN => n1603_port);
   NEXT_REGISTERS_reg_25_60_inst : DLH_X1 port map( G => n12108, D => N2685, Q 
                           => NEXT_REGISTERS_25_60_port);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => N466, CK => CLK, Q => 
                           n10155, QN => n1604_port);
   NEXT_REGISTERS_reg_25_59_inst : DLH_X1 port map( G => n12108, D => N2684, Q 
                           => NEXT_REGISTERS_25_59_port);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => N465, CK => CLK, Q => 
                           n10154, QN => n1605_port);
   NEXT_REGISTERS_reg_25_58_inst : DLH_X1 port map( G => n12108, D => N2683, Q 
                           => NEXT_REGISTERS_25_58_port);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => N464, CK => CLK, Q => 
                           n10153, QN => n1606_port);
   NEXT_REGISTERS_reg_25_57_inst : DLH_X1 port map( G => n12108, D => N2682, Q 
                           => NEXT_REGISTERS_25_57_port);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => N463, CK => CLK, Q => 
                           n10152, QN => n1607_port);
   NEXT_REGISTERS_reg_25_56_inst : DLH_X1 port map( G => n12108, D => N2681, Q 
                           => NEXT_REGISTERS_25_56_port);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => N462, CK => CLK, Q => 
                           n10151, QN => n1608_port);
   NEXT_REGISTERS_reg_25_55_inst : DLH_X1 port map( G => n12108, D => N2680, Q 
                           => NEXT_REGISTERS_25_55_port);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => N461, CK => CLK, Q => 
                           n10150, QN => n1609_port);
   NEXT_REGISTERS_reg_25_54_inst : DLH_X1 port map( G => n12108, D => N2679, Q 
                           => NEXT_REGISTERS_25_54_port);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => N460, CK => CLK, Q => 
                           n10149, QN => n1610_port);
   NEXT_REGISTERS_reg_25_53_inst : DLH_X1 port map( G => n12108, D => N2678, Q 
                           => NEXT_REGISTERS_25_53_port);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => N459, CK => CLK, Q => 
                           n10148, QN => n1611_port);
   NEXT_REGISTERS_reg_25_52_inst : DLH_X1 port map( G => n12109, D => N2677, Q 
                           => NEXT_REGISTERS_25_52_port);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => N458, CK => CLK, Q => 
                           n10147, QN => n1612_port);
   NEXT_REGISTERS_reg_25_51_inst : DLH_X1 port map( G => n12109, D => N2676, Q 
                           => NEXT_REGISTERS_25_51_port);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => N457, CK => CLK, Q => 
                           n10146, QN => n1613_port);
   NEXT_REGISTERS_reg_25_50_inst : DLH_X1 port map( G => n12109, D => N2675, Q 
                           => NEXT_REGISTERS_25_50_port);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => N456, CK => CLK, Q => 
                           n10145, QN => n1614_port);
   NEXT_REGISTERS_reg_25_49_inst : DLH_X1 port map( G => n12109, D => N2674, Q 
                           => NEXT_REGISTERS_25_49_port);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => N455, CK => CLK, Q => 
                           n10144, QN => n1615_port);
   NEXT_REGISTERS_reg_25_48_inst : DLH_X1 port map( G => n12109, D => N2673, Q 
                           => NEXT_REGISTERS_25_48_port);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => N454, CK => CLK, Q => 
                           n10143, QN => n1616_port);
   NEXT_REGISTERS_reg_25_47_inst : DLH_X1 port map( G => n12109, D => N2672, Q 
                           => NEXT_REGISTERS_25_47_port);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => N453, CK => CLK, Q => 
                           n10142, QN => n1617_port);
   NEXT_REGISTERS_reg_25_46_inst : DLH_X1 port map( G => n12109, D => N2671, Q 
                           => NEXT_REGISTERS_25_46_port);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => N452, CK => CLK, Q => 
                           n10141, QN => n1618_port);
   NEXT_REGISTERS_reg_25_45_inst : DLH_X1 port map( G => n12109, D => N2670, Q 
                           => NEXT_REGISTERS_25_45_port);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => N451, CK => CLK, Q => 
                           n10140, QN => n1619_port);
   NEXT_REGISTERS_reg_25_44_inst : DLH_X1 port map( G => n12109, D => N2669, Q 
                           => NEXT_REGISTERS_25_44_port);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => N450, CK => CLK, Q => 
                           n10139, QN => n1620_port);
   NEXT_REGISTERS_reg_25_43_inst : DLH_X1 port map( G => n12109, D => N2668, Q 
                           => NEXT_REGISTERS_25_43_port);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => N449, CK => CLK, Q => 
                           n10138, QN => n1621_port);
   NEXT_REGISTERS_reg_25_42_inst : DLH_X1 port map( G => n12109, D => N2667, Q 
                           => NEXT_REGISTERS_25_42_port);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => N448, CK => CLK, Q => 
                           n10137, QN => n1622_port);
   NEXT_REGISTERS_reg_25_41_inst : DLH_X1 port map( G => n12110, D => N2666, Q 
                           => NEXT_REGISTERS_25_41_port);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => N447, CK => CLK, Q => 
                           n10136, QN => n1623_port);
   NEXT_REGISTERS_reg_25_40_inst : DLH_X1 port map( G => n12110, D => N2665, Q 
                           => NEXT_REGISTERS_25_40_port);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => N446, CK => CLK, Q => 
                           n10135, QN => n1624_port);
   NEXT_REGISTERS_reg_25_39_inst : DLH_X1 port map( G => n12110, D => N2664, Q 
                           => NEXT_REGISTERS_25_39_port);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => N445, CK => CLK, Q => 
                           n10134, QN => n1625_port);
   NEXT_REGISTERS_reg_25_38_inst : DLH_X1 port map( G => n12110, D => N2663, Q 
                           => NEXT_REGISTERS_25_38_port);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => N444, CK => CLK, Q => 
                           n10133, QN => n1626_port);
   NEXT_REGISTERS_reg_25_37_inst : DLH_X1 port map( G => n12110, D => N2662, Q 
                           => NEXT_REGISTERS_25_37_port);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => N443, CK => CLK, Q => 
                           n10132, QN => n1627_port);
   NEXT_REGISTERS_reg_25_36_inst : DLH_X1 port map( G => n12110, D => N2661, Q 
                           => NEXT_REGISTERS_25_36_port);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => N442, CK => CLK, Q => 
                           n10131, QN => n1628_port);
   NEXT_REGISTERS_reg_25_35_inst : DLH_X1 port map( G => n12110, D => N2660, Q 
                           => NEXT_REGISTERS_25_35_port);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => N441, CK => CLK, Q => 
                           n10130, QN => n1629_port);
   NEXT_REGISTERS_reg_25_34_inst : DLH_X1 port map( G => n12110, D => N2659, Q 
                           => NEXT_REGISTERS_25_34_port);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => N440, CK => CLK, Q => 
                           n10129, QN => n1630_port);
   NEXT_REGISTERS_reg_25_33_inst : DLH_X1 port map( G => n12110, D => N2658, Q 
                           => NEXT_REGISTERS_25_33_port);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => N439, CK => CLK, Q => 
                           n10128, QN => n1631_port);
   NEXT_REGISTERS_reg_25_32_inst : DLH_X1 port map( G => n12110, D => N2657, Q 
                           => NEXT_REGISTERS_25_32_port);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => N438, CK => CLK, Q => 
                           n10127, QN => n1632_port);
   NEXT_REGISTERS_reg_25_31_inst : DLH_X1 port map( G => n12110, D => N2656, Q 
                           => NEXT_REGISTERS_25_31_port);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => N437, CK => CLK, Q => 
                           n10126, QN => n1633_port);
   NEXT_REGISTERS_reg_25_30_inst : DLH_X1 port map( G => n12111, D => N2655, Q 
                           => NEXT_REGISTERS_25_30_port);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => N436, CK => CLK, Q => 
                           n10125, QN => n1634_port);
   NEXT_REGISTERS_reg_25_29_inst : DLH_X1 port map( G => n12111, D => N2654, Q 
                           => NEXT_REGISTERS_25_29_port);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => N435, CK => CLK, Q => 
                           n10124, QN => n1635_port);
   NEXT_REGISTERS_reg_25_28_inst : DLH_X1 port map( G => n12111, D => N2653, Q 
                           => NEXT_REGISTERS_25_28_port);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => N434, CK => CLK, Q => 
                           n10123, QN => n1636_port);
   NEXT_REGISTERS_reg_25_27_inst : DLH_X1 port map( G => n12111, D => N2652, Q 
                           => NEXT_REGISTERS_25_27_port);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => N433, CK => CLK, Q => 
                           n10122, QN => n1637_port);
   NEXT_REGISTERS_reg_25_26_inst : DLH_X1 port map( G => n12111, D => N2651, Q 
                           => NEXT_REGISTERS_25_26_port);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => N432, CK => CLK, Q => 
                           n10121, QN => n1638_port);
   NEXT_REGISTERS_reg_25_25_inst : DLH_X1 port map( G => n12111, D => N2650, Q 
                           => NEXT_REGISTERS_25_25_port);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => N431, CK => CLK, Q => 
                           n10120, QN => n1639_port);
   NEXT_REGISTERS_reg_25_24_inst : DLH_X1 port map( G => n12111, D => N2649, Q 
                           => NEXT_REGISTERS_25_24_port);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => N430, CK => CLK, Q => 
                           n10119, QN => n1640_port);
   NEXT_REGISTERS_reg_25_23_inst : DLH_X1 port map( G => n12111, D => N2648, Q 
                           => NEXT_REGISTERS_25_23_port);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => N429, CK => CLK, Q => 
                           n10118, QN => n1641_port);
   NEXT_REGISTERS_reg_25_22_inst : DLH_X1 port map( G => n12111, D => N2647, Q 
                           => NEXT_REGISTERS_25_22_port);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => N428, CK => CLK, Q => 
                           n10117, QN => n1642_port);
   NEXT_REGISTERS_reg_25_21_inst : DLH_X1 port map( G => n12111, D => N2646, Q 
                           => NEXT_REGISTERS_25_21_port);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => N427, CK => CLK, Q => 
                           n10116, QN => n1643_port);
   NEXT_REGISTERS_reg_25_20_inst : DLH_X1 port map( G => n12111, D => N2645, Q 
                           => NEXT_REGISTERS_25_20_port);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => N426, CK => CLK, Q => 
                           n10115, QN => n1644_port);
   NEXT_REGISTERS_reg_25_19_inst : DLH_X1 port map( G => n12112, D => N2644, Q 
                           => NEXT_REGISTERS_25_19_port);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => N425, CK => CLK, Q => 
                           n10114, QN => n1645_port);
   NEXT_REGISTERS_reg_25_18_inst : DLH_X1 port map( G => n12112, D => N2643, Q 
                           => NEXT_REGISTERS_25_18_port);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => N424, CK => CLK, Q => 
                           n10113, QN => n1646_port);
   NEXT_REGISTERS_reg_25_17_inst : DLH_X1 port map( G => n12112, D => N2642, Q 
                           => NEXT_REGISTERS_25_17_port);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => N423, CK => CLK, Q => 
                           n10112, QN => n1647_port);
   NEXT_REGISTERS_reg_25_16_inst : DLH_X1 port map( G => n12112, D => N2641, Q 
                           => NEXT_REGISTERS_25_16_port);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => N422, CK => CLK, Q => 
                           n10111, QN => n1648_port);
   NEXT_REGISTERS_reg_25_15_inst : DLH_X1 port map( G => n12112, D => N2640, Q 
                           => NEXT_REGISTERS_25_15_port);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => N421, CK => CLK, Q => 
                           n10110, QN => n1649_port);
   NEXT_REGISTERS_reg_25_14_inst : DLH_X1 port map( G => n12112, D => N2639, Q 
                           => NEXT_REGISTERS_25_14_port);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => N420, CK => CLK, Q => 
                           n10109, QN => n1650_port);
   NEXT_REGISTERS_reg_25_13_inst : DLH_X1 port map( G => n12112, D => N2638, Q 
                           => NEXT_REGISTERS_25_13_port);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => N419, CK => CLK, Q => 
                           n10108, QN => n1651_port);
   NEXT_REGISTERS_reg_25_12_inst : DLH_X1 port map( G => n12112, D => N2637, Q 
                           => NEXT_REGISTERS_25_12_port);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => N418, CK => CLK, Q => 
                           n10107, QN => n1652_port);
   NEXT_REGISTERS_reg_25_11_inst : DLH_X1 port map( G => n12112, D => N2636, Q 
                           => NEXT_REGISTERS_25_11_port);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => N417, CK => CLK, Q => 
                           n10106, QN => n1653_port);
   NEXT_REGISTERS_reg_25_10_inst : DLH_X1 port map( G => n12112, D => N2635, Q 
                           => NEXT_REGISTERS_25_10_port);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => N416, CK => CLK, Q => 
                           n10105, QN => n1654_port);
   NEXT_REGISTERS_reg_25_9_inst : DLH_X1 port map( G => n12112, D => N2634, Q 
                           => NEXT_REGISTERS_25_9_port);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => N415, CK => CLK, Q => n10104
                           , QN => n1655_port);
   NEXT_REGISTERS_reg_25_8_inst : DLH_X1 port map( G => n12113, D => N2633, Q 
                           => NEXT_REGISTERS_25_8_port);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => N414, CK => CLK, Q => n10103
                           , QN => n1656_port);
   NEXT_REGISTERS_reg_25_7_inst : DLH_X1 port map( G => n12113, D => N2632, Q 
                           => NEXT_REGISTERS_25_7_port);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => N413, CK => CLK, Q => n10102
                           , QN => n1657_port);
   NEXT_REGISTERS_reg_25_6_inst : DLH_X1 port map( G => n12113, D => N2631, Q 
                           => NEXT_REGISTERS_25_6_port);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => N412, CK => CLK, Q => n10101
                           , QN => n1658_port);
   NEXT_REGISTERS_reg_25_5_inst : DLH_X1 port map( G => n12113, D => N2630, Q 
                           => NEXT_REGISTERS_25_5_port);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => N411, CK => CLK, Q => n10100
                           , QN => n1659_port);
   NEXT_REGISTERS_reg_25_4_inst : DLH_X1 port map( G => n12113, D => N2629, Q 
                           => NEXT_REGISTERS_25_4_port);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => N410, CK => CLK, Q => n10099
                           , QN => n1660_port);
   NEXT_REGISTERS_reg_25_3_inst : DLH_X1 port map( G => n12113, D => N2628, Q 
                           => NEXT_REGISTERS_25_3_port);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => N409, CK => CLK, Q => n10098
                           , QN => n1661_port);
   NEXT_REGISTERS_reg_25_2_inst : DLH_X1 port map( G => n12113, D => N2627, Q 
                           => NEXT_REGISTERS_25_2_port);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => N408, CK => CLK, Q => n10097
                           , QN => n1662_port);
   NEXT_REGISTERS_reg_25_1_inst : DLH_X1 port map( G => n12113, D => N2626, Q 
                           => NEXT_REGISTERS_25_1_port);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => N407, CK => CLK, Q => n10096
                           , QN => n1663_port);
   NEXT_REGISTERS_reg_25_0_inst : DLH_X1 port map( G => n12113, D => N2625, Q 
                           => NEXT_REGISTERS_25_0_port);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => N406, CK => CLK, Q => n10095
                           , QN => n1664_port);
   NEXT_REGISTERS_reg_26_63_inst : DLH_X1 port map( G => n12117, D => N2623, Q 
                           => NEXT_REGISTERS_26_63_port);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => N405, CK => CLK, Q => 
                           n10606, QN => n1665_port);
   NEXT_REGISTERS_reg_26_62_inst : DLH_X1 port map( G => n12117, D => N2622, Q 
                           => NEXT_REGISTERS_26_62_port);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => N404, CK => CLK, Q => 
                           n10605, QN => n1666_port);
   NEXT_REGISTERS_reg_26_61_inst : DLH_X1 port map( G => n12117, D => N2621, Q 
                           => NEXT_REGISTERS_26_61_port);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => N403, CK => CLK, Q => 
                           n10604, QN => n1667_port);
   NEXT_REGISTERS_reg_26_60_inst : DLH_X1 port map( G => n12117, D => N2620, Q 
                           => NEXT_REGISTERS_26_60_port);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => N402, CK => CLK, Q => 
                           n10603, QN => n1668_port);
   NEXT_REGISTERS_reg_26_59_inst : DLH_X1 port map( G => n12117, D => N2619, Q 
                           => NEXT_REGISTERS_26_59_port);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => N401, CK => CLK, Q => 
                           n10602, QN => n1669_port);
   NEXT_REGISTERS_reg_26_58_inst : DLH_X1 port map( G => n12117, D => N2618, Q 
                           => NEXT_REGISTERS_26_58_port);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => N400, CK => CLK, Q => 
                           n10601, QN => n1670_port);
   NEXT_REGISTERS_reg_26_57_inst : DLH_X1 port map( G => n12117, D => N2617, Q 
                           => NEXT_REGISTERS_26_57_port);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => N399, CK => CLK, Q => 
                           n10600, QN => n1671_port);
   NEXT_REGISTERS_reg_26_56_inst : DLH_X1 port map( G => n12117, D => N2616, Q 
                           => NEXT_REGISTERS_26_56_port);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => N398, CK => CLK, Q => 
                           n10599, QN => n1672_port);
   NEXT_REGISTERS_reg_26_55_inst : DLH_X1 port map( G => n12117, D => N2615, Q 
                           => NEXT_REGISTERS_26_55_port);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => N397, CK => CLK, Q => 
                           n10598, QN => n1673_port);
   NEXT_REGISTERS_reg_26_54_inst : DLH_X1 port map( G => n12117, D => N2614, Q 
                           => NEXT_REGISTERS_26_54_port);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => N396, CK => CLK, Q => 
                           n10597, QN => n1674_port);
   NEXT_REGISTERS_reg_26_53_inst : DLH_X1 port map( G => n12117, D => N2613, Q 
                           => NEXT_REGISTERS_26_53_port);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => N395, CK => CLK, Q => 
                           n10596, QN => n1675_port);
   NEXT_REGISTERS_reg_26_52_inst : DLH_X1 port map( G => n12118, D => N2612, Q 
                           => NEXT_REGISTERS_26_52_port);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => N394, CK => CLK, Q => 
                           n10595, QN => n1676_port);
   NEXT_REGISTERS_reg_26_51_inst : DLH_X1 port map( G => n12118, D => N2611, Q 
                           => NEXT_REGISTERS_26_51_port);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => N393, CK => CLK, Q => 
                           n10594, QN => n1677_port);
   NEXT_REGISTERS_reg_26_50_inst : DLH_X1 port map( G => n12118, D => N2610, Q 
                           => NEXT_REGISTERS_26_50_port);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => N392, CK => CLK, Q => 
                           n10593, QN => n1678_port);
   NEXT_REGISTERS_reg_26_49_inst : DLH_X1 port map( G => n12118, D => N2609, Q 
                           => NEXT_REGISTERS_26_49_port);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => N391, CK => CLK, Q => 
                           n10592, QN => n1679_port);
   NEXT_REGISTERS_reg_26_48_inst : DLH_X1 port map( G => n12118, D => N2608, Q 
                           => NEXT_REGISTERS_26_48_port);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => N390, CK => CLK, Q => 
                           n10591, QN => n1680_port);
   NEXT_REGISTERS_reg_26_47_inst : DLH_X1 port map( G => n12118, D => N2607, Q 
                           => NEXT_REGISTERS_26_47_port);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => N389, CK => CLK, Q => 
                           n10590, QN => n1681_port);
   NEXT_REGISTERS_reg_26_46_inst : DLH_X1 port map( G => n12118, D => N2606, Q 
                           => NEXT_REGISTERS_26_46_port);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => N388, CK => CLK, Q => 
                           n10589, QN => n1682_port);
   NEXT_REGISTERS_reg_26_45_inst : DLH_X1 port map( G => n12118, D => N2605, Q 
                           => NEXT_REGISTERS_26_45_port);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => N387, CK => CLK, Q => 
                           n10588, QN => n1683_port);
   NEXT_REGISTERS_reg_26_44_inst : DLH_X1 port map( G => n12118, D => N2604, Q 
                           => NEXT_REGISTERS_26_44_port);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => N386, CK => CLK, Q => 
                           n10587, QN => n1684_port);
   NEXT_REGISTERS_reg_26_43_inst : DLH_X1 port map( G => n12118, D => N2603, Q 
                           => NEXT_REGISTERS_26_43_port);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => N385, CK => CLK, Q => 
                           n10586, QN => n1685_port);
   NEXT_REGISTERS_reg_26_42_inst : DLH_X1 port map( G => n12118, D => N2602, Q 
                           => NEXT_REGISTERS_26_42_port);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => N384, CK => CLK, Q => 
                           n10585, QN => n1686_port);
   NEXT_REGISTERS_reg_26_41_inst : DLH_X1 port map( G => n12119, D => N2601, Q 
                           => NEXT_REGISTERS_26_41_port);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => N383, CK => CLK, Q => 
                           n10584, QN => n1687_port);
   NEXT_REGISTERS_reg_26_40_inst : DLH_X1 port map( G => n12119, D => N2600, Q 
                           => NEXT_REGISTERS_26_40_port);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => N382, CK => CLK, Q => 
                           n10583, QN => n1688_port);
   NEXT_REGISTERS_reg_26_39_inst : DLH_X1 port map( G => n12119, D => N2599, Q 
                           => NEXT_REGISTERS_26_39_port);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => N381, CK => CLK, Q => 
                           n10582, QN => n1689_port);
   NEXT_REGISTERS_reg_26_38_inst : DLH_X1 port map( G => n12119, D => N2598, Q 
                           => NEXT_REGISTERS_26_38_port);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => N380, CK => CLK, Q => 
                           n10581, QN => n1690_port);
   NEXT_REGISTERS_reg_26_37_inst : DLH_X1 port map( G => n12119, D => N2597, Q 
                           => NEXT_REGISTERS_26_37_port);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => N379, CK => CLK, Q => 
                           n10580, QN => n1691_port);
   NEXT_REGISTERS_reg_26_36_inst : DLH_X1 port map( G => n12119, D => N2596, Q 
                           => NEXT_REGISTERS_26_36_port);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => N378, CK => CLK, Q => 
                           n10579, QN => n1692_port);
   NEXT_REGISTERS_reg_26_35_inst : DLH_X1 port map( G => n12119, D => N2595, Q 
                           => NEXT_REGISTERS_26_35_port);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => N377, CK => CLK, Q => 
                           n10578, QN => n1693_port);
   NEXT_REGISTERS_reg_26_34_inst : DLH_X1 port map( G => n12119, D => N2594, Q 
                           => NEXT_REGISTERS_26_34_port);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => N376, CK => CLK, Q => 
                           n10577, QN => n1694_port);
   NEXT_REGISTERS_reg_26_33_inst : DLH_X1 port map( G => n12119, D => N2593, Q 
                           => NEXT_REGISTERS_26_33_port);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => N375, CK => CLK, Q => 
                           n10576, QN => n1695_port);
   NEXT_REGISTERS_reg_26_32_inst : DLH_X1 port map( G => n12119, D => N2592, Q 
                           => NEXT_REGISTERS_26_32_port);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => N374, CK => CLK, Q => 
                           n10575, QN => n1696_port);
   NEXT_REGISTERS_reg_26_31_inst : DLH_X1 port map( G => n12119, D => N2591, Q 
                           => NEXT_REGISTERS_26_31_port);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => N373, CK => CLK, Q => 
                           n10574, QN => n1697_port);
   NEXT_REGISTERS_reg_26_30_inst : DLH_X1 port map( G => n12120, D => N2590, Q 
                           => NEXT_REGISTERS_26_30_port);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => N372, CK => CLK, Q => 
                           n10573, QN => n1698_port);
   NEXT_REGISTERS_reg_26_29_inst : DLH_X1 port map( G => n12120, D => N2589, Q 
                           => NEXT_REGISTERS_26_29_port);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => N371, CK => CLK, Q => 
                           n10572, QN => n1699_port);
   NEXT_REGISTERS_reg_26_28_inst : DLH_X1 port map( G => n12120, D => N2588, Q 
                           => NEXT_REGISTERS_26_28_port);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => N370, CK => CLK, Q => 
                           n10571, QN => n1700_port);
   NEXT_REGISTERS_reg_26_27_inst : DLH_X1 port map( G => n12120, D => N2587, Q 
                           => NEXT_REGISTERS_26_27_port);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => N369, CK => CLK, Q => 
                           n10570, QN => n1701_port);
   NEXT_REGISTERS_reg_26_26_inst : DLH_X1 port map( G => n12120, D => N2586, Q 
                           => NEXT_REGISTERS_26_26_port);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => N368, CK => CLK, Q => 
                           n10569, QN => n1702_port);
   NEXT_REGISTERS_reg_26_25_inst : DLH_X1 port map( G => n12120, D => N2585, Q 
                           => NEXT_REGISTERS_26_25_port);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => N367, CK => CLK, Q => 
                           n10568, QN => n1703_port);
   NEXT_REGISTERS_reg_26_24_inst : DLH_X1 port map( G => n12120, D => N2584, Q 
                           => NEXT_REGISTERS_26_24_port);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => N366, CK => CLK, Q => 
                           n10567, QN => n1704_port);
   NEXT_REGISTERS_reg_26_23_inst : DLH_X1 port map( G => n12120, D => N2583, Q 
                           => NEXT_REGISTERS_26_23_port);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => N365, CK => CLK, Q => 
                           n10566, QN => n1705_port);
   NEXT_REGISTERS_reg_26_22_inst : DLH_X1 port map( G => n12120, D => N2582, Q 
                           => NEXT_REGISTERS_26_22_port);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => N364, CK => CLK, Q => 
                           n10565, QN => n1706_port);
   NEXT_REGISTERS_reg_26_21_inst : DLH_X1 port map( G => n12120, D => N2581, Q 
                           => NEXT_REGISTERS_26_21_port);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => N363, CK => CLK, Q => 
                           n10564, QN => n1707_port);
   NEXT_REGISTERS_reg_26_20_inst : DLH_X1 port map( G => n12120, D => N2580, Q 
                           => NEXT_REGISTERS_26_20_port);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => N362, CK => CLK, Q => 
                           n10563, QN => n1708_port);
   NEXT_REGISTERS_reg_26_19_inst : DLH_X1 port map( G => n12121, D => N2579, Q 
                           => NEXT_REGISTERS_26_19_port);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => N361, CK => CLK, Q => 
                           n10562, QN => n1709_port);
   NEXT_REGISTERS_reg_26_18_inst : DLH_X1 port map( G => n12121, D => N2578, Q 
                           => NEXT_REGISTERS_26_18_port);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => N360, CK => CLK, Q => 
                           n10561, QN => n1710_port);
   NEXT_REGISTERS_reg_26_17_inst : DLH_X1 port map( G => n12121, D => N2577, Q 
                           => NEXT_REGISTERS_26_17_port);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => N359, CK => CLK, Q => 
                           n10560, QN => n1711_port);
   NEXT_REGISTERS_reg_26_16_inst : DLH_X1 port map( G => n12121, D => N2576, Q 
                           => NEXT_REGISTERS_26_16_port);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => N358, CK => CLK, Q => 
                           n10559, QN => n1712_port);
   NEXT_REGISTERS_reg_26_15_inst : DLH_X1 port map( G => n12121, D => N2575, Q 
                           => NEXT_REGISTERS_26_15_port);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => N357, CK => CLK, Q => 
                           n10558, QN => n1713_port);
   NEXT_REGISTERS_reg_26_14_inst : DLH_X1 port map( G => n12121, D => N2574, Q 
                           => NEXT_REGISTERS_26_14_port);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => N356, CK => CLK, Q => 
                           n10557, QN => n1714_port);
   NEXT_REGISTERS_reg_26_13_inst : DLH_X1 port map( G => n12121, D => N2573, Q 
                           => NEXT_REGISTERS_26_13_port);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => N355, CK => CLK, Q => 
                           n10556, QN => n1715_port);
   NEXT_REGISTERS_reg_26_12_inst : DLH_X1 port map( G => n12121, D => N2572, Q 
                           => NEXT_REGISTERS_26_12_port);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => N354, CK => CLK, Q => 
                           n10555, QN => n1716_port);
   NEXT_REGISTERS_reg_26_11_inst : DLH_X1 port map( G => n12121, D => N2571, Q 
                           => NEXT_REGISTERS_26_11_port);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => N353, CK => CLK, Q => 
                           n10554, QN => n1717_port);
   NEXT_REGISTERS_reg_26_10_inst : DLH_X1 port map( G => n12121, D => N2570, Q 
                           => NEXT_REGISTERS_26_10_port);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => N352, CK => CLK, Q => 
                           n10553, QN => n1718_port);
   NEXT_REGISTERS_reg_26_9_inst : DLH_X1 port map( G => n12121, D => N2569, Q 
                           => NEXT_REGISTERS_26_9_port);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => N351, CK => CLK, Q => n10552
                           , QN => n1719_port);
   NEXT_REGISTERS_reg_26_8_inst : DLH_X1 port map( G => n12122, D => N2568, Q 
                           => NEXT_REGISTERS_26_8_port);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => N350, CK => CLK, Q => n10551
                           , QN => n1720_port);
   NEXT_REGISTERS_reg_26_7_inst : DLH_X1 port map( G => n12122, D => N2567, Q 
                           => NEXT_REGISTERS_26_7_port);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => N349, CK => CLK, Q => n10550
                           , QN => n1721_port);
   NEXT_REGISTERS_reg_26_6_inst : DLH_X1 port map( G => n12122, D => N2566, Q 
                           => NEXT_REGISTERS_26_6_port);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => N348, CK => CLK, Q => n10549
                           , QN => n1722_port);
   NEXT_REGISTERS_reg_26_5_inst : DLH_X1 port map( G => n12122, D => N2565, Q 
                           => NEXT_REGISTERS_26_5_port);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => N347, CK => CLK, Q => n10548
                           , QN => n1723_port);
   NEXT_REGISTERS_reg_26_4_inst : DLH_X1 port map( G => n12122, D => N2564, Q 
                           => NEXT_REGISTERS_26_4_port);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => N346, CK => CLK, Q => n10547
                           , QN => n1724_port);
   NEXT_REGISTERS_reg_26_3_inst : DLH_X1 port map( G => n12122, D => N2563, Q 
                           => NEXT_REGISTERS_26_3_port);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => N345, CK => CLK, Q => n10546
                           , QN => n1725_port);
   NEXT_REGISTERS_reg_26_2_inst : DLH_X1 port map( G => n12122, D => N2562, Q 
                           => NEXT_REGISTERS_26_2_port);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => N344, CK => CLK, Q => n10545
                           , QN => n1726_port);
   NEXT_REGISTERS_reg_26_1_inst : DLH_X1 port map( G => n12122, D => N2561, Q 
                           => NEXT_REGISTERS_26_1_port);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => N343, CK => CLK, Q => n10544
                           , QN => n1727_port);
   NEXT_REGISTERS_reg_26_0_inst : DLH_X1 port map( G => n12122, D => N2560, Q 
                           => NEXT_REGISTERS_26_0_port);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => N342, CK => CLK, Q => n10543
                           , QN => n1728_port);
   NEXT_REGISTERS_reg_27_63_inst : DLH_X1 port map( G => n12126, D => N2558, Q 
                           => NEXT_REGISTERS_27_63_port);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => N341, CK => CLK, Q => n9710
                           , QN => n1729_port);
   NEXT_REGISTERS_reg_27_62_inst : DLH_X1 port map( G => n12126, D => N2557, Q 
                           => NEXT_REGISTERS_27_62_port);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => N340, CK => CLK, Q => n9709
                           , QN => n1730_port);
   NEXT_REGISTERS_reg_27_61_inst : DLH_X1 port map( G => n12126, D => N2556, Q 
                           => NEXT_REGISTERS_27_61_port);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => N339, CK => CLK, Q => n9708
                           , QN => n1731_port);
   NEXT_REGISTERS_reg_27_60_inst : DLH_X1 port map( G => n12126, D => N2555, Q 
                           => NEXT_REGISTERS_27_60_port);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => N338, CK => CLK, Q => n9707
                           , QN => n1732_port);
   NEXT_REGISTERS_reg_27_59_inst : DLH_X1 port map( G => n12126, D => N2554, Q 
                           => NEXT_REGISTERS_27_59_port);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => N337, CK => CLK, Q => n9706
                           , QN => n1733_port);
   NEXT_REGISTERS_reg_27_58_inst : DLH_X1 port map( G => n12126, D => N2553, Q 
                           => NEXT_REGISTERS_27_58_port);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => N336, CK => CLK, Q => n9705
                           , QN => n1734_port);
   NEXT_REGISTERS_reg_27_57_inst : DLH_X1 port map( G => n12126, D => N2552, Q 
                           => NEXT_REGISTERS_27_57_port);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => N335, CK => CLK, Q => n9704
                           , QN => n1735_port);
   NEXT_REGISTERS_reg_27_56_inst : DLH_X1 port map( G => n12126, D => N2551, Q 
                           => NEXT_REGISTERS_27_56_port);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => N334, CK => CLK, Q => n9703
                           , QN => n1736_port);
   NEXT_REGISTERS_reg_27_55_inst : DLH_X1 port map( G => n12126, D => N2550, Q 
                           => NEXT_REGISTERS_27_55_port);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => N333, CK => CLK, Q => n9702
                           , QN => n1737_port);
   NEXT_REGISTERS_reg_27_54_inst : DLH_X1 port map( G => n12126, D => N2549, Q 
                           => NEXT_REGISTERS_27_54_port);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => N332, CK => CLK, Q => n9701
                           , QN => n1738_port);
   NEXT_REGISTERS_reg_27_53_inst : DLH_X1 port map( G => n12126, D => N2548, Q 
                           => NEXT_REGISTERS_27_53_port);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => N331, CK => CLK, Q => n9700
                           , QN => n1739_port);
   NEXT_REGISTERS_reg_27_52_inst : DLH_X1 port map( G => n12127, D => N2547, Q 
                           => NEXT_REGISTERS_27_52_port);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => N330, CK => CLK, Q => n9699
                           , QN => n1740_port);
   NEXT_REGISTERS_reg_27_51_inst : DLH_X1 port map( G => n12127, D => N2546, Q 
                           => NEXT_REGISTERS_27_51_port);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => N329, CK => CLK, Q => n9698
                           , QN => n1741_port);
   NEXT_REGISTERS_reg_27_50_inst : DLH_X1 port map( G => n12127, D => N2545, Q 
                           => NEXT_REGISTERS_27_50_port);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => N328, CK => CLK, Q => n9697
                           , QN => n1742_port);
   NEXT_REGISTERS_reg_27_49_inst : DLH_X1 port map( G => n12127, D => N2544, Q 
                           => NEXT_REGISTERS_27_49_port);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => N327, CK => CLK, Q => n9696
                           , QN => n1743_port);
   NEXT_REGISTERS_reg_27_48_inst : DLH_X1 port map( G => n12127, D => N2543, Q 
                           => NEXT_REGISTERS_27_48_port);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => N326, CK => CLK, Q => n9695
                           , QN => n1744_port);
   NEXT_REGISTERS_reg_27_47_inst : DLH_X1 port map( G => n12127, D => N2542, Q 
                           => NEXT_REGISTERS_27_47_port);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => N325, CK => CLK, Q => n9694
                           , QN => n1745_port);
   NEXT_REGISTERS_reg_27_46_inst : DLH_X1 port map( G => n12127, D => N2541, Q 
                           => NEXT_REGISTERS_27_46_port);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => N324, CK => CLK, Q => n9693
                           , QN => n1746_port);
   NEXT_REGISTERS_reg_27_45_inst : DLH_X1 port map( G => n12127, D => N2540, Q 
                           => NEXT_REGISTERS_27_45_port);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => N323, CK => CLK, Q => n9692
                           , QN => n1747_port);
   NEXT_REGISTERS_reg_27_44_inst : DLH_X1 port map( G => n12127, D => N2539, Q 
                           => NEXT_REGISTERS_27_44_port);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => N322, CK => CLK, Q => n9691
                           , QN => n1748_port);
   NEXT_REGISTERS_reg_27_43_inst : DLH_X1 port map( G => n12127, D => N2538, Q 
                           => NEXT_REGISTERS_27_43_port);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => N321, CK => CLK, Q => n9690
                           , QN => n1749_port);
   NEXT_REGISTERS_reg_27_42_inst : DLH_X1 port map( G => n12127, D => N2537, Q 
                           => NEXT_REGISTERS_27_42_port);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => N320, CK => CLK, Q => n9689
                           , QN => n1750_port);
   NEXT_REGISTERS_reg_27_41_inst : DLH_X1 port map( G => n12128, D => N2536, Q 
                           => NEXT_REGISTERS_27_41_port);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => N319, CK => CLK, Q => n9688
                           , QN => n1751_port);
   NEXT_REGISTERS_reg_27_40_inst : DLH_X1 port map( G => n12128, D => N2535, Q 
                           => NEXT_REGISTERS_27_40_port);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => N318, CK => CLK, Q => n9687
                           , QN => n1752_port);
   NEXT_REGISTERS_reg_27_39_inst : DLH_X1 port map( G => n12128, D => N2534, Q 
                           => NEXT_REGISTERS_27_39_port);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => N317, CK => CLK, Q => n9686
                           , QN => n1753_port);
   NEXT_REGISTERS_reg_27_38_inst : DLH_X1 port map( G => n12128, D => N2533, Q 
                           => NEXT_REGISTERS_27_38_port);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => N316, CK => CLK, Q => n9685
                           , QN => n1754_port);
   NEXT_REGISTERS_reg_27_37_inst : DLH_X1 port map( G => n12128, D => N2532, Q 
                           => NEXT_REGISTERS_27_37_port);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => N315, CK => CLK, Q => n9684
                           , QN => n1755_port);
   NEXT_REGISTERS_reg_27_36_inst : DLH_X1 port map( G => n12128, D => N2531, Q 
                           => NEXT_REGISTERS_27_36_port);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => N314, CK => CLK, Q => n9683
                           , QN => n1756_port);
   NEXT_REGISTERS_reg_27_35_inst : DLH_X1 port map( G => n12128, D => N2530, Q 
                           => NEXT_REGISTERS_27_35_port);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => N313, CK => CLK, Q => n9682
                           , QN => n1757_port);
   NEXT_REGISTERS_reg_27_34_inst : DLH_X1 port map( G => n12128, D => N2529, Q 
                           => NEXT_REGISTERS_27_34_port);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => N312, CK => CLK, Q => n9681
                           , QN => n1758_port);
   NEXT_REGISTERS_reg_27_33_inst : DLH_X1 port map( G => n12128, D => N2528, Q 
                           => NEXT_REGISTERS_27_33_port);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => N311, CK => CLK, Q => n9680
                           , QN => n1759_port);
   NEXT_REGISTERS_reg_27_32_inst : DLH_X1 port map( G => n12128, D => N2527, Q 
                           => NEXT_REGISTERS_27_32_port);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => N310, CK => CLK, Q => n9679
                           , QN => n1760_port);
   NEXT_REGISTERS_reg_27_31_inst : DLH_X1 port map( G => n12128, D => N2526, Q 
                           => NEXT_REGISTERS_27_31_port);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => N309, CK => CLK, Q => n9678
                           , QN => n1761_port);
   NEXT_REGISTERS_reg_27_30_inst : DLH_X1 port map( G => n12129, D => N2525, Q 
                           => NEXT_REGISTERS_27_30_port);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => N308, CK => CLK, Q => n9677
                           , QN => n1762_port);
   NEXT_REGISTERS_reg_27_29_inst : DLH_X1 port map( G => n12129, D => N2524, Q 
                           => NEXT_REGISTERS_27_29_port);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => N307, CK => CLK, Q => n9676
                           , QN => n1763_port);
   NEXT_REGISTERS_reg_27_28_inst : DLH_X1 port map( G => n12129, D => N2523, Q 
                           => NEXT_REGISTERS_27_28_port);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => N306, CK => CLK, Q => n9675
                           , QN => n1764_port);
   NEXT_REGISTERS_reg_27_27_inst : DLH_X1 port map( G => n12129, D => N2522, Q 
                           => NEXT_REGISTERS_27_27_port);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => N305, CK => CLK, Q => n9674
                           , QN => n1765_port);
   NEXT_REGISTERS_reg_27_26_inst : DLH_X1 port map( G => n12129, D => N2521, Q 
                           => NEXT_REGISTERS_27_26_port);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => N304, CK => CLK, Q => n9673
                           , QN => n1766_port);
   NEXT_REGISTERS_reg_27_25_inst : DLH_X1 port map( G => n12129, D => N2520, Q 
                           => NEXT_REGISTERS_27_25_port);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => N303, CK => CLK, Q => n9672
                           , QN => n1767_port);
   NEXT_REGISTERS_reg_27_24_inst : DLH_X1 port map( G => n12129, D => N2519, Q 
                           => NEXT_REGISTERS_27_24_port);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => N302, CK => CLK, Q => n9671
                           , QN => n1768_port);
   NEXT_REGISTERS_reg_27_23_inst : DLH_X1 port map( G => n12129, D => N2518, Q 
                           => NEXT_REGISTERS_27_23_port);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => N301, CK => CLK, Q => n9670
                           , QN => n1769_port);
   NEXT_REGISTERS_reg_27_22_inst : DLH_X1 port map( G => n12129, D => N2517, Q 
                           => NEXT_REGISTERS_27_22_port);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => N300, CK => CLK, Q => n9669
                           , QN => n1770_port);
   NEXT_REGISTERS_reg_27_21_inst : DLH_X1 port map( G => n12129, D => N2516, Q 
                           => NEXT_REGISTERS_27_21_port);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => N299, CK => CLK, Q => n9668
                           , QN => n1771_port);
   NEXT_REGISTERS_reg_27_20_inst : DLH_X1 port map( G => n12129, D => N2515, Q 
                           => NEXT_REGISTERS_27_20_port);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => N298, CK => CLK, Q => n9667
                           , QN => n1772_port);
   NEXT_REGISTERS_reg_27_19_inst : DLH_X1 port map( G => n12130, D => N2514, Q 
                           => NEXT_REGISTERS_27_19_port);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => N297, CK => CLK, Q => n9666
                           , QN => n1773_port);
   NEXT_REGISTERS_reg_27_18_inst : DLH_X1 port map( G => n12130, D => N2513, Q 
                           => NEXT_REGISTERS_27_18_port);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => N296, CK => CLK, Q => n9665
                           , QN => n1774_port);
   NEXT_REGISTERS_reg_27_17_inst : DLH_X1 port map( G => n12130, D => N2512, Q 
                           => NEXT_REGISTERS_27_17_port);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => N295, CK => CLK, Q => n9664
                           , QN => n1775_port);
   NEXT_REGISTERS_reg_27_16_inst : DLH_X1 port map( G => n12130, D => N2511, Q 
                           => NEXT_REGISTERS_27_16_port);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => N294, CK => CLK, Q => n9663
                           , QN => n1776_port);
   NEXT_REGISTERS_reg_27_15_inst : DLH_X1 port map( G => n12130, D => N2510, Q 
                           => NEXT_REGISTERS_27_15_port);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => N293, CK => CLK, Q => n9662
                           , QN => n1777_port);
   NEXT_REGISTERS_reg_27_14_inst : DLH_X1 port map( G => n12130, D => N2509, Q 
                           => NEXT_REGISTERS_27_14_port);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => N292, CK => CLK, Q => n9661
                           , QN => n1778_port);
   NEXT_REGISTERS_reg_27_13_inst : DLH_X1 port map( G => n12130, D => N2508, Q 
                           => NEXT_REGISTERS_27_13_port);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => N291, CK => CLK, Q => n9660
                           , QN => n1779_port);
   NEXT_REGISTERS_reg_27_12_inst : DLH_X1 port map( G => n12130, D => N2507, Q 
                           => NEXT_REGISTERS_27_12_port);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => N290, CK => CLK, Q => n9659
                           , QN => n1780_port);
   NEXT_REGISTERS_reg_27_11_inst : DLH_X1 port map( G => n12130, D => N2506, Q 
                           => NEXT_REGISTERS_27_11_port);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => N289, CK => CLK, Q => n9658
                           , QN => n1781_port);
   NEXT_REGISTERS_reg_27_10_inst : DLH_X1 port map( G => n12130, D => N2505, Q 
                           => NEXT_REGISTERS_27_10_port);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => N288, CK => CLK, Q => n9657
                           , QN => n1782_port);
   NEXT_REGISTERS_reg_27_9_inst : DLH_X1 port map( G => n12130, D => N2504, Q 
                           => NEXT_REGISTERS_27_9_port);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => N287, CK => CLK, Q => n9656,
                           QN => n1783_port);
   NEXT_REGISTERS_reg_27_8_inst : DLH_X1 port map( G => n12131, D => N2503, Q 
                           => NEXT_REGISTERS_27_8_port);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => N286, CK => CLK, Q => n9655,
                           QN => n1784_port);
   NEXT_REGISTERS_reg_27_7_inst : DLH_X1 port map( G => n12131, D => N2502, Q 
                           => NEXT_REGISTERS_27_7_port);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => N285, CK => CLK, Q => n9654,
                           QN => n1785_port);
   NEXT_REGISTERS_reg_27_6_inst : DLH_X1 port map( G => n12131, D => N2501, Q 
                           => NEXT_REGISTERS_27_6_port);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => N284, CK => CLK, Q => n9653,
                           QN => n1786_port);
   NEXT_REGISTERS_reg_27_5_inst : DLH_X1 port map( G => n12131, D => N2500, Q 
                           => NEXT_REGISTERS_27_5_port);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => N283, CK => CLK, Q => n9652,
                           QN => n1787_port);
   NEXT_REGISTERS_reg_27_4_inst : DLH_X1 port map( G => n12131, D => N2499, Q 
                           => NEXT_REGISTERS_27_4_port);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => N282, CK => CLK, Q => n9651,
                           QN => n1788_port);
   NEXT_REGISTERS_reg_27_3_inst : DLH_X1 port map( G => n12131, D => N2498, Q 
                           => NEXT_REGISTERS_27_3_port);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => N281, CK => CLK, Q => n9650,
                           QN => n1789_port);
   NEXT_REGISTERS_reg_27_2_inst : DLH_X1 port map( G => n12131, D => N2497, Q 
                           => NEXT_REGISTERS_27_2_port);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => N280, CK => CLK, Q => n9649,
                           QN => n1790_port);
   NEXT_REGISTERS_reg_27_1_inst : DLH_X1 port map( G => n12131, D => N2496, Q 
                           => NEXT_REGISTERS_27_1_port);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => N279, CK => CLK, Q => n9648,
                           QN => n1791_port);
   NEXT_REGISTERS_reg_27_0_inst : DLH_X1 port map( G => n12131, D => N2495, Q 
                           => NEXT_REGISTERS_27_0_port);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => N278, CK => CLK, Q => n9647,
                           QN => n1792_port);
   NEXT_REGISTERS_reg_28_63_inst : DLH_X1 port map( G => n12135, D => N2493, Q 
                           => NEXT_REGISTERS_28_63_port);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => N277, CK => CLK, Q => 
                           n_1832, QN => n1793_port);
   NEXT_REGISTERS_reg_28_62_inst : DLH_X1 port map( G => n12135, D => N2492, Q 
                           => NEXT_REGISTERS_28_62_port);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => N276, CK => CLK, Q => 
                           n_1833, QN => n1794_port);
   NEXT_REGISTERS_reg_28_61_inst : DLH_X1 port map( G => n12135, D => N2491, Q 
                           => NEXT_REGISTERS_28_61_port);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => N275, CK => CLK, Q => 
                           n_1834, QN => n1795_port);
   NEXT_REGISTERS_reg_28_60_inst : DLH_X1 port map( G => n12135, D => N2490, Q 
                           => NEXT_REGISTERS_28_60_port);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => N274, CK => CLK, Q => 
                           n_1835, QN => n1796_port);
   NEXT_REGISTERS_reg_28_59_inst : DLH_X1 port map( G => n12135, D => N2489, Q 
                           => NEXT_REGISTERS_28_59_port);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => N273, CK => CLK, Q => 
                           n_1836, QN => n1797_port);
   NEXT_REGISTERS_reg_28_58_inst : DLH_X1 port map( G => n12135, D => N2488, Q 
                           => NEXT_REGISTERS_28_58_port);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => N272, CK => CLK, Q => 
                           n_1837, QN => n1798_port);
   NEXT_REGISTERS_reg_28_57_inst : DLH_X1 port map( G => n12135, D => N2487, Q 
                           => NEXT_REGISTERS_28_57_port);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => N271, CK => CLK, Q => 
                           n_1838, QN => n1799_port);
   NEXT_REGISTERS_reg_28_56_inst : DLH_X1 port map( G => n12135, D => N2486, Q 
                           => NEXT_REGISTERS_28_56_port);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => N270, CK => CLK, Q => 
                           n_1839, QN => n1800_port);
   NEXT_REGISTERS_reg_28_55_inst : DLH_X1 port map( G => n12135, D => N2485, Q 
                           => NEXT_REGISTERS_28_55_port);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => N269, CK => CLK, Q => 
                           n_1840, QN => n1801_port);
   NEXT_REGISTERS_reg_28_54_inst : DLH_X1 port map( G => n12135, D => N2484, Q 
                           => NEXT_REGISTERS_28_54_port);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => N268, CK => CLK, Q => 
                           n_1841, QN => n1802_port);
   NEXT_REGISTERS_reg_28_53_inst : DLH_X1 port map( G => n12135, D => N2483, Q 
                           => NEXT_REGISTERS_28_53_port);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => N267, CK => CLK, Q => 
                           n_1842, QN => n1803_port);
   NEXT_REGISTERS_reg_28_52_inst : DLH_X1 port map( G => n12136, D => N2482, Q 
                           => NEXT_REGISTERS_28_52_port);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => N266, CK => CLK, Q => 
                           n_1843, QN => n1804_port);
   NEXT_REGISTERS_reg_28_51_inst : DLH_X1 port map( G => n12136, D => N2481, Q 
                           => NEXT_REGISTERS_28_51_port);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => N265, CK => CLK, Q => 
                           n_1844, QN => n1805_port);
   NEXT_REGISTERS_reg_28_50_inst : DLH_X1 port map( G => n12136, D => N2480, Q 
                           => NEXT_REGISTERS_28_50_port);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => N264, CK => CLK, Q => 
                           n_1845, QN => n1806_port);
   NEXT_REGISTERS_reg_28_49_inst : DLH_X1 port map( G => n12136, D => N2479, Q 
                           => NEXT_REGISTERS_28_49_port);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => N263, CK => CLK, Q => 
                           n_1846, QN => n1807_port);
   NEXT_REGISTERS_reg_28_48_inst : DLH_X1 port map( G => n12136, D => N2478, Q 
                           => NEXT_REGISTERS_28_48_port);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => N262, CK => CLK, Q => 
                           n_1847, QN => n1808_port);
   NEXT_REGISTERS_reg_28_47_inst : DLH_X1 port map( G => n12136, D => N2477, Q 
                           => NEXT_REGISTERS_28_47_port);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => N261, CK => CLK, Q => 
                           n_1848, QN => n1809_port);
   NEXT_REGISTERS_reg_28_46_inst : DLH_X1 port map( G => n12136, D => N2476, Q 
                           => NEXT_REGISTERS_28_46_port);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => N260, CK => CLK, Q => 
                           n_1849, QN => n1810_port);
   NEXT_REGISTERS_reg_28_45_inst : DLH_X1 port map( G => n12136, D => N2475, Q 
                           => NEXT_REGISTERS_28_45_port);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => N259, CK => CLK, Q => 
                           n_1850, QN => n1811_port);
   NEXT_REGISTERS_reg_28_44_inst : DLH_X1 port map( G => n12136, D => N2474, Q 
                           => NEXT_REGISTERS_28_44_port);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => N258, CK => CLK, Q => 
                           n_1851, QN => n1812_port);
   NEXT_REGISTERS_reg_28_43_inst : DLH_X1 port map( G => n12136, D => N2473, Q 
                           => NEXT_REGISTERS_28_43_port);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => N257, CK => CLK, Q => 
                           n_1852, QN => n1813_port);
   NEXT_REGISTERS_reg_28_42_inst : DLH_X1 port map( G => n12136, D => N2472, Q 
                           => NEXT_REGISTERS_28_42_port);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => N256, CK => CLK, Q => 
                           n_1853, QN => n1814_port);
   NEXT_REGISTERS_reg_28_41_inst : DLH_X1 port map( G => n12137, D => N2471, Q 
                           => NEXT_REGISTERS_28_41_port);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => N255, CK => CLK, Q => 
                           n_1854, QN => n1815_port);
   NEXT_REGISTERS_reg_28_40_inst : DLH_X1 port map( G => n12137, D => N2470, Q 
                           => NEXT_REGISTERS_28_40_port);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => N254, CK => CLK, Q => 
                           n_1855, QN => n1816_port);
   NEXT_REGISTERS_reg_28_39_inst : DLH_X1 port map( G => n12137, D => N2469, Q 
                           => NEXT_REGISTERS_28_39_port);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => N253, CK => CLK, Q => 
                           n_1856, QN => n1817_port);
   NEXT_REGISTERS_reg_28_38_inst : DLH_X1 port map( G => n12137, D => N2468, Q 
                           => NEXT_REGISTERS_28_38_port);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => N252, CK => CLK, Q => 
                           n_1857, QN => n1818_port);
   NEXT_REGISTERS_reg_28_37_inst : DLH_X1 port map( G => n12137, D => N2467, Q 
                           => NEXT_REGISTERS_28_37_port);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => N251, CK => CLK, Q => 
                           n_1858, QN => n1819_port);
   NEXT_REGISTERS_reg_28_36_inst : DLH_X1 port map( G => n12137, D => N2466, Q 
                           => NEXT_REGISTERS_28_36_port);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => N250, CK => CLK, Q => 
                           n_1859, QN => n1820_port);
   NEXT_REGISTERS_reg_28_35_inst : DLH_X1 port map( G => n12137, D => N2465, Q 
                           => NEXT_REGISTERS_28_35_port);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => N249, CK => CLK, Q => 
                           n_1860, QN => n1821_port);
   NEXT_REGISTERS_reg_28_34_inst : DLH_X1 port map( G => n12137, D => N2464, Q 
                           => NEXT_REGISTERS_28_34_port);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => N248, CK => CLK, Q => 
                           n_1861, QN => n1822_port);
   NEXT_REGISTERS_reg_28_33_inst : DLH_X1 port map( G => n12137, D => N2463, Q 
                           => NEXT_REGISTERS_28_33_port);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => N247, CK => CLK, Q => 
                           n_1862, QN => n1823_port);
   NEXT_REGISTERS_reg_28_32_inst : DLH_X1 port map( G => n12137, D => N2462, Q 
                           => NEXT_REGISTERS_28_32_port);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => N246, CK => CLK, Q => 
                           n_1863, QN => n1824_port);
   NEXT_REGISTERS_reg_28_31_inst : DLH_X1 port map( G => n12137, D => N2461, Q 
                           => NEXT_REGISTERS_28_31_port);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => N245, CK => CLK, Q => 
                           n_1864, QN => n1825_port);
   NEXT_REGISTERS_reg_28_30_inst : DLH_X1 port map( G => n12138, D => N2460, Q 
                           => NEXT_REGISTERS_28_30_port);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => N244, CK => CLK, Q => 
                           n_1865, QN => n1826_port);
   NEXT_REGISTERS_reg_28_29_inst : DLH_X1 port map( G => n12138, D => N2459, Q 
                           => NEXT_REGISTERS_28_29_port);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => N243, CK => CLK, Q => 
                           n_1866, QN => n1827_port);
   NEXT_REGISTERS_reg_28_28_inst : DLH_X1 port map( G => n12138, D => N2458, Q 
                           => NEXT_REGISTERS_28_28_port);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => N242, CK => CLK, Q => 
                           n_1867, QN => n1828_port);
   NEXT_REGISTERS_reg_28_27_inst : DLH_X1 port map( G => n12138, D => N2457, Q 
                           => NEXT_REGISTERS_28_27_port);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => N241, CK => CLK, Q => 
                           n_1868, QN => n1829_port);
   NEXT_REGISTERS_reg_28_26_inst : DLH_X1 port map( G => n12138, D => N2456, Q 
                           => NEXT_REGISTERS_28_26_port);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => N240, CK => CLK, Q => 
                           n_1869, QN => n1830_port);
   NEXT_REGISTERS_reg_28_25_inst : DLH_X1 port map( G => n12138, D => N2455, Q 
                           => NEXT_REGISTERS_28_25_port);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => N239, CK => CLK, Q => 
                           n_1870, QN => n1831_port);
   NEXT_REGISTERS_reg_28_24_inst : DLH_X1 port map( G => n12138, D => N2454, Q 
                           => NEXT_REGISTERS_28_24_port);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => N238, CK => CLK, Q => 
                           n_1871, QN => n1832_port);
   NEXT_REGISTERS_reg_28_23_inst : DLH_X1 port map( G => n12138, D => N2453, Q 
                           => NEXT_REGISTERS_28_23_port);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => N237, CK => CLK, Q => 
                           n_1872, QN => n1833_port);
   NEXT_REGISTERS_reg_28_22_inst : DLH_X1 port map( G => n12138, D => N2452, Q 
                           => NEXT_REGISTERS_28_22_port);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => N236, CK => CLK, Q => 
                           n_1873, QN => n1834_port);
   NEXT_REGISTERS_reg_28_21_inst : DLH_X1 port map( G => n12138, D => N2451, Q 
                           => NEXT_REGISTERS_28_21_port);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => N235, CK => CLK, Q => 
                           n_1874, QN => n1835_port);
   NEXT_REGISTERS_reg_28_20_inst : DLH_X1 port map( G => n12138, D => N2450, Q 
                           => NEXT_REGISTERS_28_20_port);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => N234, CK => CLK, Q => 
                           n_1875, QN => n1836_port);
   NEXT_REGISTERS_reg_28_19_inst : DLH_X1 port map( G => n12139, D => N2449, Q 
                           => NEXT_REGISTERS_28_19_port);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => N233, CK => CLK, Q => 
                           n_1876, QN => n1837_port);
   NEXT_REGISTERS_reg_28_18_inst : DLH_X1 port map( G => n12139, D => N2448, Q 
                           => NEXT_REGISTERS_28_18_port);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => N232, CK => CLK, Q => 
                           n_1877, QN => n1838_port);
   NEXT_REGISTERS_reg_28_17_inst : DLH_X1 port map( G => n12139, D => N2447, Q 
                           => NEXT_REGISTERS_28_17_port);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => N231, CK => CLK, Q => 
                           n_1878, QN => n1839_port);
   NEXT_REGISTERS_reg_28_16_inst : DLH_X1 port map( G => n12139, D => N2446, Q 
                           => NEXT_REGISTERS_28_16_port);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => N230, CK => CLK, Q => 
                           n_1879, QN => n1840_port);
   NEXT_REGISTERS_reg_28_15_inst : DLH_X1 port map( G => n12139, D => N2445, Q 
                           => NEXT_REGISTERS_28_15_port);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => N229, CK => CLK, Q => 
                           n_1880, QN => n1841_port);
   NEXT_REGISTERS_reg_28_14_inst : DLH_X1 port map( G => n12139, D => N2444, Q 
                           => NEXT_REGISTERS_28_14_port);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => N228, CK => CLK, Q => 
                           n_1881, QN => n1842_port);
   NEXT_REGISTERS_reg_28_13_inst : DLH_X1 port map( G => n12139, D => N2443, Q 
                           => NEXT_REGISTERS_28_13_port);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => N227, CK => CLK, Q => 
                           n_1882, QN => n1843_port);
   NEXT_REGISTERS_reg_28_12_inst : DLH_X1 port map( G => n12139, D => N2442, Q 
                           => NEXT_REGISTERS_28_12_port);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => N226, CK => CLK, Q => 
                           n_1883, QN => n1844_port);
   NEXT_REGISTERS_reg_28_11_inst : DLH_X1 port map( G => n12139, D => N2441, Q 
                           => NEXT_REGISTERS_28_11_port);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => N225, CK => CLK, Q => 
                           n_1884, QN => n1845_port);
   NEXT_REGISTERS_reg_28_10_inst : DLH_X1 port map( G => n12139, D => N2440, Q 
                           => NEXT_REGISTERS_28_10_port);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => N224, CK => CLK, Q => 
                           n_1885, QN => n1846_port);
   NEXT_REGISTERS_reg_28_9_inst : DLH_X1 port map( G => n12139, D => N2439, Q 
                           => NEXT_REGISTERS_28_9_port);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => N223, CK => CLK, Q => n_1886
                           , QN => n1847_port);
   NEXT_REGISTERS_reg_28_8_inst : DLH_X1 port map( G => n12140, D => N2438, Q 
                           => NEXT_REGISTERS_28_8_port);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => N222, CK => CLK, Q => n_1887
                           , QN => n1848_port);
   NEXT_REGISTERS_reg_28_7_inst : DLH_X1 port map( G => n12140, D => N2437, Q 
                           => NEXT_REGISTERS_28_7_port);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => N221, CK => CLK, Q => n_1888
                           , QN => n1849_port);
   NEXT_REGISTERS_reg_28_6_inst : DLH_X1 port map( G => n12140, D => N2436, Q 
                           => NEXT_REGISTERS_28_6_port);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => N220, CK => CLK, Q => n_1889
                           , QN => n1850_port);
   NEXT_REGISTERS_reg_28_5_inst : DLH_X1 port map( G => n12140, D => N2435, Q 
                           => NEXT_REGISTERS_28_5_port);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => N219, CK => CLK, Q => n_1890
                           , QN => n1851_port);
   NEXT_REGISTERS_reg_28_4_inst : DLH_X1 port map( G => n12140, D => N2434, Q 
                           => NEXT_REGISTERS_28_4_port);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => N218, CK => CLK, Q => n_1891
                           , QN => n1852_port);
   NEXT_REGISTERS_reg_28_3_inst : DLH_X1 port map( G => n12140, D => N2433, Q 
                           => NEXT_REGISTERS_28_3_port);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => N217, CK => CLK, Q => n_1892
                           , QN => n1853_port);
   NEXT_REGISTERS_reg_28_2_inst : DLH_X1 port map( G => n12140, D => N2432, Q 
                           => NEXT_REGISTERS_28_2_port);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => N216, CK => CLK, Q => n_1893
                           , QN => n1854_port);
   NEXT_REGISTERS_reg_28_1_inst : DLH_X1 port map( G => n12140, D => N2431, Q 
                           => NEXT_REGISTERS_28_1_port);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => N215, CK => CLK, Q => n_1894
                           , QN => n1855_port);
   NEXT_REGISTERS_reg_28_0_inst : DLH_X1 port map( G => n12140, D => N2430, Q 
                           => NEXT_REGISTERS_28_0_port);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => N214, CK => CLK, Q => n_1895
                           , QN => n1856_port);
   NEXT_REGISTERS_reg_29_63_inst : DLH_X1 port map( G => n12144, D => N2428, Q 
                           => NEXT_REGISTERS_29_63_port);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => N213, CK => CLK, Q => 
                           n_1896, QN => n1857_port);
   NEXT_REGISTERS_reg_29_62_inst : DLH_X1 port map( G => n12144, D => N2427, Q 
                           => NEXT_REGISTERS_29_62_port);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => N212, CK => CLK, Q => 
                           n_1897, QN => n1858_port);
   NEXT_REGISTERS_reg_29_61_inst : DLH_X1 port map( G => n12144, D => N2426, Q 
                           => NEXT_REGISTERS_29_61_port);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => N211, CK => CLK, Q => 
                           n_1898, QN => n1859_port);
   NEXT_REGISTERS_reg_29_60_inst : DLH_X1 port map( G => n12144, D => N2425, Q 
                           => NEXT_REGISTERS_29_60_port);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => N210, CK => CLK, Q => 
                           n_1899, QN => n1860_port);
   NEXT_REGISTERS_reg_29_59_inst : DLH_X1 port map( G => n12144, D => N2424, Q 
                           => NEXT_REGISTERS_29_59_port);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => N209, CK => CLK, Q => 
                           n_1900, QN => n1861_port);
   NEXT_REGISTERS_reg_29_58_inst : DLH_X1 port map( G => n12144, D => N2423, Q 
                           => NEXT_REGISTERS_29_58_port);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => N208, CK => CLK, Q => 
                           n_1901, QN => n1862_port);
   NEXT_REGISTERS_reg_29_57_inst : DLH_X1 port map( G => n12144, D => N2422, Q 
                           => NEXT_REGISTERS_29_57_port);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => N207, CK => CLK, Q => 
                           n_1902, QN => n1863_port);
   NEXT_REGISTERS_reg_29_56_inst : DLH_X1 port map( G => n12144, D => N2421, Q 
                           => NEXT_REGISTERS_29_56_port);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => N206, CK => CLK, Q => 
                           n_1903, QN => n1864_port);
   NEXT_REGISTERS_reg_29_55_inst : DLH_X1 port map( G => n12144, D => N2420, Q 
                           => NEXT_REGISTERS_29_55_port);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => N205, CK => CLK, Q => 
                           n_1904, QN => n1865_port);
   NEXT_REGISTERS_reg_29_54_inst : DLH_X1 port map( G => n12144, D => N2419, Q 
                           => NEXT_REGISTERS_29_54_port);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => N204, CK => CLK, Q => 
                           n_1905, QN => n1866_port);
   NEXT_REGISTERS_reg_29_53_inst : DLH_X1 port map( G => n12144, D => N2418, Q 
                           => NEXT_REGISTERS_29_53_port);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => N203, CK => CLK, Q => 
                           n_1906, QN => n1867_port);
   NEXT_REGISTERS_reg_29_52_inst : DLH_X1 port map( G => n12145, D => N2417, Q 
                           => NEXT_REGISTERS_29_52_port);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => N202, CK => CLK, Q => 
                           n_1907, QN => n1868_port);
   NEXT_REGISTERS_reg_29_51_inst : DLH_X1 port map( G => n12145, D => N2416, Q 
                           => NEXT_REGISTERS_29_51_port);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => N201, CK => CLK, Q => 
                           n_1908, QN => n1869_port);
   NEXT_REGISTERS_reg_29_50_inst : DLH_X1 port map( G => n12145, D => N2415, Q 
                           => NEXT_REGISTERS_29_50_port);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => N200, CK => CLK, Q => 
                           n_1909, QN => n1870_port);
   NEXT_REGISTERS_reg_29_49_inst : DLH_X1 port map( G => n12145, D => N2414, Q 
                           => NEXT_REGISTERS_29_49_port);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => N199, CK => CLK, Q => 
                           n_1910, QN => n1871_port);
   NEXT_REGISTERS_reg_29_48_inst : DLH_X1 port map( G => n12145, D => N2413, Q 
                           => NEXT_REGISTERS_29_48_port);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => N198, CK => CLK, Q => 
                           n_1911, QN => n1872_port);
   NEXT_REGISTERS_reg_29_47_inst : DLH_X1 port map( G => n12145, D => N2412, Q 
                           => NEXT_REGISTERS_29_47_port);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => N197, CK => CLK, Q => 
                           n_1912, QN => n1873_port);
   NEXT_REGISTERS_reg_29_46_inst : DLH_X1 port map( G => n12145, D => N2411, Q 
                           => NEXT_REGISTERS_29_46_port);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => N196, CK => CLK, Q => 
                           n_1913, QN => n1874_port);
   NEXT_REGISTERS_reg_29_45_inst : DLH_X1 port map( G => n12145, D => N2410, Q 
                           => NEXT_REGISTERS_29_45_port);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => N195, CK => CLK, Q => 
                           n_1914, QN => n1875_port);
   NEXT_REGISTERS_reg_29_44_inst : DLH_X1 port map( G => n12145, D => N2409, Q 
                           => NEXT_REGISTERS_29_44_port);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => N194, CK => CLK, Q => 
                           n_1915, QN => n1876_port);
   NEXT_REGISTERS_reg_29_43_inst : DLH_X1 port map( G => n12145, D => N2408, Q 
                           => NEXT_REGISTERS_29_43_port);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => N193, CK => CLK, Q => 
                           n_1916, QN => n1877_port);
   NEXT_REGISTERS_reg_29_42_inst : DLH_X1 port map( G => n12145, D => N2407, Q 
                           => NEXT_REGISTERS_29_42_port);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => N192, CK => CLK, Q => 
                           n_1917, QN => n1878_port);
   NEXT_REGISTERS_reg_29_41_inst : DLH_X1 port map( G => n12146, D => N2406, Q 
                           => NEXT_REGISTERS_29_41_port);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => N191, CK => CLK, Q => 
                           n_1918, QN => n1879_port);
   NEXT_REGISTERS_reg_29_40_inst : DLH_X1 port map( G => n12146, D => N2405, Q 
                           => NEXT_REGISTERS_29_40_port);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => N190, CK => CLK, Q => 
                           n_1919, QN => n1880_port);
   NEXT_REGISTERS_reg_29_39_inst : DLH_X1 port map( G => n12146, D => N2404, Q 
                           => NEXT_REGISTERS_29_39_port);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => N189, CK => CLK, Q => 
                           n_1920, QN => n1881_port);
   NEXT_REGISTERS_reg_29_38_inst : DLH_X1 port map( G => n12146, D => N2403, Q 
                           => NEXT_REGISTERS_29_38_port);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => N188, CK => CLK, Q => 
                           n_1921, QN => n1882_port);
   NEXT_REGISTERS_reg_29_37_inst : DLH_X1 port map( G => n12146, D => N2402, Q 
                           => NEXT_REGISTERS_29_37_port);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => N187, CK => CLK, Q => 
                           n_1922, QN => n1883_port);
   NEXT_REGISTERS_reg_29_36_inst : DLH_X1 port map( G => n12146, D => N2401, Q 
                           => NEXT_REGISTERS_29_36_port);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => N186, CK => CLK, Q => 
                           n_1923, QN => n1884_port);
   NEXT_REGISTERS_reg_29_35_inst : DLH_X1 port map( G => n12146, D => N2400, Q 
                           => NEXT_REGISTERS_29_35_port);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => N185, CK => CLK, Q => 
                           n_1924, QN => n1885_port);
   NEXT_REGISTERS_reg_29_34_inst : DLH_X1 port map( G => n12146, D => N2399, Q 
                           => NEXT_REGISTERS_29_34_port);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => N184, CK => CLK, Q => 
                           n_1925, QN => n1886_port);
   NEXT_REGISTERS_reg_29_33_inst : DLH_X1 port map( G => n12146, D => N2398, Q 
                           => NEXT_REGISTERS_29_33_port);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => N183, CK => CLK, Q => 
                           n_1926, QN => n1887_port);
   NEXT_REGISTERS_reg_29_32_inst : DLH_X1 port map( G => n12146, D => N2397, Q 
                           => NEXT_REGISTERS_29_32_port);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => N182, CK => CLK, Q => 
                           n_1927, QN => n1888_port);
   NEXT_REGISTERS_reg_29_31_inst : DLH_X1 port map( G => n12146, D => N2396, Q 
                           => NEXT_REGISTERS_29_31_port);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => N181, CK => CLK, Q => 
                           n_1928, QN => n1889_port);
   NEXT_REGISTERS_reg_29_30_inst : DLH_X1 port map( G => n12147, D => N2395, Q 
                           => NEXT_REGISTERS_29_30_port);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => N180, CK => CLK, Q => 
                           n_1929, QN => n1890_port);
   NEXT_REGISTERS_reg_29_29_inst : DLH_X1 port map( G => n12147, D => N2394, Q 
                           => NEXT_REGISTERS_29_29_port);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => N179, CK => CLK, Q => 
                           n_1930, QN => n1891_port);
   NEXT_REGISTERS_reg_29_28_inst : DLH_X1 port map( G => n12147, D => N2393, Q 
                           => NEXT_REGISTERS_29_28_port);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => N178, CK => CLK, Q => 
                           n_1931, QN => n1892_port);
   NEXT_REGISTERS_reg_29_27_inst : DLH_X1 port map( G => n12147, D => N2392, Q 
                           => NEXT_REGISTERS_29_27_port);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => N177, CK => CLK, Q => 
                           n_1932, QN => n1893_port);
   NEXT_REGISTERS_reg_29_26_inst : DLH_X1 port map( G => n12147, D => N2391, Q 
                           => NEXT_REGISTERS_29_26_port);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => N176, CK => CLK, Q => 
                           n_1933, QN => n1894_port);
   NEXT_REGISTERS_reg_29_25_inst : DLH_X1 port map( G => n12147, D => N2390, Q 
                           => NEXT_REGISTERS_29_25_port);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => N175, CK => CLK, Q => 
                           n_1934, QN => n1895_port);
   NEXT_REGISTERS_reg_29_24_inst : DLH_X1 port map( G => n12147, D => N2389, Q 
                           => NEXT_REGISTERS_29_24_port);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => N174, CK => CLK, Q => 
                           n_1935, QN => n1896_port);
   NEXT_REGISTERS_reg_29_23_inst : DLH_X1 port map( G => n12147, D => N2388, Q 
                           => NEXT_REGISTERS_29_23_port);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => N173, CK => CLK, Q => 
                           n_1936, QN => n1897_port);
   NEXT_REGISTERS_reg_29_22_inst : DLH_X1 port map( G => n12147, D => N2387, Q 
                           => NEXT_REGISTERS_29_22_port);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => N172, CK => CLK, Q => 
                           n_1937, QN => n1898_port);
   NEXT_REGISTERS_reg_29_21_inst : DLH_X1 port map( G => n12147, D => N2386, Q 
                           => NEXT_REGISTERS_29_21_port);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => N171, CK => CLK, Q => 
                           n_1938, QN => n1899_port);
   NEXT_REGISTERS_reg_29_20_inst : DLH_X1 port map( G => n12147, D => N2385, Q 
                           => NEXT_REGISTERS_29_20_port);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => N170, CK => CLK, Q => 
                           n_1939, QN => n1900_port);
   NEXT_REGISTERS_reg_29_19_inst : DLH_X1 port map( G => n12148, D => N2384, Q 
                           => NEXT_REGISTERS_29_19_port);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => N169, CK => CLK, Q => 
                           n_1940, QN => n1901_port);
   NEXT_REGISTERS_reg_29_18_inst : DLH_X1 port map( G => n12148, D => N2383, Q 
                           => NEXT_REGISTERS_29_18_port);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => N168, CK => CLK, Q => 
                           n_1941, QN => n1902_port);
   NEXT_REGISTERS_reg_29_17_inst : DLH_X1 port map( G => n12148, D => N2382, Q 
                           => NEXT_REGISTERS_29_17_port);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => N167, CK => CLK, Q => 
                           n_1942, QN => n1903_port);
   NEXT_REGISTERS_reg_29_16_inst : DLH_X1 port map( G => n12148, D => N2381, Q 
                           => NEXT_REGISTERS_29_16_port);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => N166, CK => CLK, Q => 
                           n_1943, QN => n1904_port);
   NEXT_REGISTERS_reg_29_15_inst : DLH_X1 port map( G => n12148, D => N2380, Q 
                           => NEXT_REGISTERS_29_15_port);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => N165, CK => CLK, Q => 
                           n_1944, QN => n1905_port);
   NEXT_REGISTERS_reg_29_14_inst : DLH_X1 port map( G => n12148, D => N2379, Q 
                           => NEXT_REGISTERS_29_14_port);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => N164, CK => CLK, Q => 
                           n_1945, QN => n1906_port);
   NEXT_REGISTERS_reg_29_13_inst : DLH_X1 port map( G => n12148, D => N2378, Q 
                           => NEXT_REGISTERS_29_13_port);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => N163, CK => CLK, Q => 
                           n_1946, QN => n1907_port);
   NEXT_REGISTERS_reg_29_12_inst : DLH_X1 port map( G => n12148, D => N2377, Q 
                           => NEXT_REGISTERS_29_12_port);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => N162, CK => CLK, Q => 
                           n_1947, QN => n1908_port);
   NEXT_REGISTERS_reg_29_11_inst : DLH_X1 port map( G => n12148, D => N2376, Q 
                           => NEXT_REGISTERS_29_11_port);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => N161, CK => CLK, Q => 
                           n_1948, QN => n1909_port);
   NEXT_REGISTERS_reg_29_10_inst : DLH_X1 port map( G => n12148, D => N2375, Q 
                           => NEXT_REGISTERS_29_10_port);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => N160, CK => CLK, Q => 
                           n_1949, QN => n1910_port);
   NEXT_REGISTERS_reg_29_9_inst : DLH_X1 port map( G => n12148, D => N2374, Q 
                           => NEXT_REGISTERS_29_9_port);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => N159, CK => CLK, Q => n_1950
                           , QN => n1911_port);
   NEXT_REGISTERS_reg_29_8_inst : DLH_X1 port map( G => n12149, D => N2373, Q 
                           => NEXT_REGISTERS_29_8_port);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => N158, CK => CLK, Q => n_1951
                           , QN => n1912_port);
   NEXT_REGISTERS_reg_29_7_inst : DLH_X1 port map( G => n12149, D => N2372, Q 
                           => NEXT_REGISTERS_29_7_port);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => N157, CK => CLK, Q => n_1952
                           , QN => n1913_port);
   NEXT_REGISTERS_reg_29_6_inst : DLH_X1 port map( G => n12149, D => N2371, Q 
                           => NEXT_REGISTERS_29_6_port);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => N156, CK => CLK, Q => n_1953
                           , QN => n1914_port);
   NEXT_REGISTERS_reg_29_5_inst : DLH_X1 port map( G => n12149, D => N2370, Q 
                           => NEXT_REGISTERS_29_5_port);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => N155, CK => CLK, Q => n_1954
                           , QN => n1915_port);
   NEXT_REGISTERS_reg_29_4_inst : DLH_X1 port map( G => n12149, D => N2369, Q 
                           => NEXT_REGISTERS_29_4_port);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => N154, CK => CLK, Q => n_1955
                           , QN => n1916_port);
   NEXT_REGISTERS_reg_29_3_inst : DLH_X1 port map( G => n12149, D => N2368, Q 
                           => NEXT_REGISTERS_29_3_port);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => N153, CK => CLK, Q => n_1956
                           , QN => n1917_port);
   NEXT_REGISTERS_reg_29_2_inst : DLH_X1 port map( G => n12149, D => N2367, Q 
                           => NEXT_REGISTERS_29_2_port);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => N152, CK => CLK, Q => n_1957
                           , QN => n1918_port);
   NEXT_REGISTERS_reg_29_1_inst : DLH_X1 port map( G => n12149, D => N2366, Q 
                           => NEXT_REGISTERS_29_1_port);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => N151, CK => CLK, Q => n_1958
                           , QN => n1919_port);
   NEXT_REGISTERS_reg_29_0_inst : DLH_X1 port map( G => n12149, D => N2365, Q 
                           => NEXT_REGISTERS_29_0_port);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => N150, CK => CLK, Q => n_1959
                           , QN => n1920_port);
   NEXT_REGISTERS_reg_30_63_inst : DLH_X1 port map( G => n12158, D => N2363, Q 
                           => NEXT_REGISTERS_30_63_port);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => N149, CK => CLK, Q => 
                           n_1960, QN => n1921_port);
   NEXT_REGISTERS_reg_30_62_inst : DLH_X1 port map( G => n12158, D => N2362, Q 
                           => NEXT_REGISTERS_30_62_port);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => N148, CK => CLK, Q => 
                           n_1961, QN => n1922_port);
   NEXT_REGISTERS_reg_30_61_inst : DLH_X1 port map( G => n12158, D => N2361, Q 
                           => NEXT_REGISTERS_30_61_port);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => N147, CK => CLK, Q => 
                           n_1962, QN => n1923_port);
   NEXT_REGISTERS_reg_30_60_inst : DLH_X1 port map( G => n12158, D => N2360, Q 
                           => NEXT_REGISTERS_30_60_port);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => N146, CK => CLK, Q => 
                           n_1963, QN => n1924_port);
   NEXT_REGISTERS_reg_30_59_inst : DLH_X1 port map( G => n12158, D => N2359, Q 
                           => NEXT_REGISTERS_30_59_port);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => N145, CK => CLK, Q => 
                           n_1964, QN => n1925_port);
   NEXT_REGISTERS_reg_30_58_inst : DLH_X1 port map( G => n12158, D => N2358, Q 
                           => NEXT_REGISTERS_30_58_port);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => N144, CK => CLK, Q => 
                           n_1965, QN => n1926_port);
   NEXT_REGISTERS_reg_30_57_inst : DLH_X1 port map( G => n12158, D => N2357, Q 
                           => NEXT_REGISTERS_30_57_port);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => N143, CK => CLK, Q => 
                           n_1966, QN => n1927_port);
   NEXT_REGISTERS_reg_30_56_inst : DLH_X1 port map( G => n12158, D => N2356, Q 
                           => NEXT_REGISTERS_30_56_port);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => N142, CK => CLK, Q => 
                           n_1967, QN => n1928_port);
   NEXT_REGISTERS_reg_30_55_inst : DLH_X1 port map( G => n12158, D => N2355, Q 
                           => NEXT_REGISTERS_30_55_port);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => N141, CK => CLK, Q => 
                           n_1968, QN => n1929_port);
   NEXT_REGISTERS_reg_30_54_inst : DLH_X1 port map( G => n12157, D => N2354, Q 
                           => NEXT_REGISTERS_30_54_port);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => N140, CK => CLK, Q => 
                           n_1969, QN => n1930_port);
   NEXT_REGISTERS_reg_30_53_inst : DLH_X1 port map( G => n12157, D => N2353, Q 
                           => NEXT_REGISTERS_30_53_port);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => N139, CK => CLK, Q => 
                           n_1970, QN => n1931_port);
   NEXT_REGISTERS_reg_30_52_inst : DLH_X1 port map( G => n12157, D => N2352, Q 
                           => NEXT_REGISTERS_30_52_port);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => N138, CK => CLK, Q => 
                           n_1971, QN => n1932_port);
   NEXT_REGISTERS_reg_30_51_inst : DLH_X1 port map( G => n12157, D => N2351, Q 
                           => NEXT_REGISTERS_30_51_port);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => N137, CK => CLK, Q => 
                           n_1972, QN => n1933_port);
   NEXT_REGISTERS_reg_30_50_inst : DLH_X1 port map( G => n12157, D => N2350, Q 
                           => NEXT_REGISTERS_30_50_port);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => N136, CK => CLK, Q => 
                           n_1973, QN => n1934_port);
   NEXT_REGISTERS_reg_30_49_inst : DLH_X1 port map( G => n12157, D => N2349, Q 
                           => NEXT_REGISTERS_30_49_port);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => N135, CK => CLK, Q => 
                           n_1974, QN => n1935_port);
   NEXT_REGISTERS_reg_30_48_inst : DLH_X1 port map( G => n12157, D => N2348, Q 
                           => NEXT_REGISTERS_30_48_port);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => N134, CK => CLK, Q => 
                           n_1975, QN => n1936_port);
   NEXT_REGISTERS_reg_30_47_inst : DLH_X1 port map( G => n12157, D => N2347, Q 
                           => NEXT_REGISTERS_30_47_port);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => N133, CK => CLK, Q => 
                           n_1976, QN => n1937_port);
   NEXT_REGISTERS_reg_30_46_inst : DLH_X1 port map( G => n12157, D => N2346, Q 
                           => NEXT_REGISTERS_30_46_port);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => N132, CK => CLK, Q => 
                           n_1977, QN => n1938_port);
   NEXT_REGISTERS_reg_30_45_inst : DLH_X1 port map( G => n12157, D => N2345, Q 
                           => NEXT_REGISTERS_30_45_port);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => N131, CK => CLK, Q => 
                           n_1978, QN => n1939_port);
   NEXT_REGISTERS_reg_30_44_inst : DLH_X1 port map( G => n12157, D => N2344, Q 
                           => NEXT_REGISTERS_30_44_port);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => N130, CK => CLK, Q => 
                           n_1979, QN => n1940_port);
   NEXT_REGISTERS_reg_30_43_inst : DLH_X1 port map( G => n12156, D => N2343, Q 
                           => NEXT_REGISTERS_30_43_port);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => N129, CK => CLK, Q => 
                           n_1980, QN => n1941_port);
   NEXT_REGISTERS_reg_30_42_inst : DLH_X1 port map( G => n12156, D => N2342, Q 
                           => NEXT_REGISTERS_30_42_port);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => N128, CK => CLK, Q => 
                           n_1981, QN => n1942_port);
   NEXT_REGISTERS_reg_30_41_inst : DLH_X1 port map( G => n12156, D => N2341, Q 
                           => NEXT_REGISTERS_30_41_port);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => N127, CK => CLK, Q => 
                           n_1982, QN => n1943_port);
   NEXT_REGISTERS_reg_30_40_inst : DLH_X1 port map( G => n12156, D => N2340, Q 
                           => NEXT_REGISTERS_30_40_port);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => N126, CK => CLK, Q => 
                           n_1983, QN => n1944_port);
   NEXT_REGISTERS_reg_30_39_inst : DLH_X1 port map( G => n12156, D => N2339, Q 
                           => NEXT_REGISTERS_30_39_port);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => N125, CK => CLK, Q => 
                           n_1984, QN => n1945_port);
   NEXT_REGISTERS_reg_30_38_inst : DLH_X1 port map( G => n12156, D => N2338, Q 
                           => NEXT_REGISTERS_30_38_port);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => N124, CK => CLK, Q => 
                           n_1985, QN => n1946_port);
   NEXT_REGISTERS_reg_30_37_inst : DLH_X1 port map( G => n12156, D => N2337, Q 
                           => NEXT_REGISTERS_30_37_port);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => N123, CK => CLK, Q => 
                           n_1986, QN => n1947_port);
   NEXT_REGISTERS_reg_30_36_inst : DLH_X1 port map( G => n12156, D => N2336, Q 
                           => NEXT_REGISTERS_30_36_port);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => N122, CK => CLK, Q => 
                           n_1987, QN => n1948_port);
   NEXT_REGISTERS_reg_30_35_inst : DLH_X1 port map( G => n12156, D => N2335, Q 
                           => NEXT_REGISTERS_30_35_port);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => N121, CK => CLK, Q => 
                           n_1988, QN => n1949_port);
   NEXT_REGISTERS_reg_30_34_inst : DLH_X1 port map( G => n12156, D => N2334, Q 
                           => NEXT_REGISTERS_30_34_port);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => N120, CK => CLK, Q => 
                           n_1989, QN => n1950_port);
   NEXT_REGISTERS_reg_30_33_inst : DLH_X1 port map( G => n12156, D => N2333, Q 
                           => NEXT_REGISTERS_30_33_port);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => N119, CK => CLK, Q => 
                           n_1990, QN => n1951_port);
   NEXT_REGISTERS_reg_30_32_inst : DLH_X1 port map( G => n12155, D => N2332, Q 
                           => NEXT_REGISTERS_30_32_port);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => N118, CK => CLK, Q => 
                           n_1991, QN => n1952_port);
   NEXT_REGISTERS_reg_30_31_inst : DLH_X1 port map( G => n12155, D => N2331, Q 
                           => NEXT_REGISTERS_30_31_port);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => N117, CK => CLK, Q => 
                           n_1992, QN => n1953_port);
   NEXT_REGISTERS_reg_30_30_inst : DLH_X1 port map( G => n12155, D => N2330, Q 
                           => NEXT_REGISTERS_30_30_port);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => N116, CK => CLK, Q => 
                           n_1993, QN => n1954_port);
   NEXT_REGISTERS_reg_30_29_inst : DLH_X1 port map( G => n12155, D => N2329, Q 
                           => NEXT_REGISTERS_30_29_port);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => N115, CK => CLK, Q => 
                           n_1994, QN => n1955_port);
   NEXT_REGISTERS_reg_30_28_inst : DLH_X1 port map( G => n12155, D => N2328, Q 
                           => NEXT_REGISTERS_30_28_port);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => N114, CK => CLK, Q => 
                           n_1995, QN => n1956_port);
   NEXT_REGISTERS_reg_30_27_inst : DLH_X1 port map( G => n12155, D => N2327, Q 
                           => NEXT_REGISTERS_30_27_port);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => N113, CK => CLK, Q => 
                           n_1996, QN => n1957_port);
   NEXT_REGISTERS_reg_30_26_inst : DLH_X1 port map( G => n12155, D => N2326, Q 
                           => NEXT_REGISTERS_30_26_port);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => N112, CK => CLK, Q => 
                           n_1997, QN => n1958_port);
   NEXT_REGISTERS_reg_30_25_inst : DLH_X1 port map( G => n12155, D => N2325, Q 
                           => NEXT_REGISTERS_30_25_port);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => N111, CK => CLK, Q => 
                           n_1998, QN => n1959_port);
   NEXT_REGISTERS_reg_30_24_inst : DLH_X1 port map( G => n12155, D => N2324, Q 
                           => NEXT_REGISTERS_30_24_port);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => N110, CK => CLK, Q => 
                           n_1999, QN => n1960_port);
   NEXT_REGISTERS_reg_30_23_inst : DLH_X1 port map( G => n12155, D => N2323, Q 
                           => NEXT_REGISTERS_30_23_port);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => N109, CK => CLK, Q => 
                           n_2000, QN => n1961_port);
   NEXT_REGISTERS_reg_30_22_inst : DLH_X1 port map( G => n12155, D => N2322, Q 
                           => NEXT_REGISTERS_30_22_port);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => N108, CK => CLK, Q => 
                           n_2001, QN => n1962_port);
   NEXT_REGISTERS_reg_30_21_inst : DLH_X1 port map( G => n12154, D => N2321, Q 
                           => NEXT_REGISTERS_30_21_port);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => N107, CK => CLK, Q => 
                           n_2002, QN => n1963_port);
   NEXT_REGISTERS_reg_30_20_inst : DLH_X1 port map( G => n12154, D => N2320, Q 
                           => NEXT_REGISTERS_30_20_port);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => N106, CK => CLK, Q => 
                           n_2003, QN => n1964_port);
   NEXT_REGISTERS_reg_30_19_inst : DLH_X1 port map( G => n12154, D => N2319, Q 
                           => NEXT_REGISTERS_30_19_port);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => N105, CK => CLK, Q => 
                           n_2004, QN => n1965_port);
   NEXT_REGISTERS_reg_30_18_inst : DLH_X1 port map( G => n12154, D => N2318, Q 
                           => NEXT_REGISTERS_30_18_port);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => N104, CK => CLK, Q => 
                           n_2005, QN => n1966_port);
   NEXT_REGISTERS_reg_30_17_inst : DLH_X1 port map( G => n12154, D => N2317, Q 
                           => NEXT_REGISTERS_30_17_port);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => N103, CK => CLK, Q => 
                           n_2006, QN => n1967_port);
   NEXT_REGISTERS_reg_30_16_inst : DLH_X1 port map( G => n12154, D => N2316, Q 
                           => NEXT_REGISTERS_30_16_port);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => N102, CK => CLK, Q => 
                           n_2007, QN => n1968_port);
   NEXT_REGISTERS_reg_30_15_inst : DLH_X1 port map( G => n12154, D => N2315, Q 
                           => NEXT_REGISTERS_30_15_port);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => N101, CK => CLK, Q => 
                           n_2008, QN => n1969_port);
   NEXT_REGISTERS_reg_30_14_inst : DLH_X1 port map( G => n12154, D => N2314, Q 
                           => NEXT_REGISTERS_30_14_port);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => N100, CK => CLK, Q => 
                           n_2009, QN => n1970_port);
   NEXT_REGISTERS_reg_30_13_inst : DLH_X1 port map( G => n12154, D => N2313, Q 
                           => NEXT_REGISTERS_30_13_port);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => N99, CK => CLK, Q => n_2010
                           , QN => n1971_port);
   NEXT_REGISTERS_reg_30_12_inst : DLH_X1 port map( G => n12154, D => N2312, Q 
                           => NEXT_REGISTERS_30_12_port);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => N98, CK => CLK, Q => n_2011
                           , QN => n1972_port);
   NEXT_REGISTERS_reg_30_11_inst : DLH_X1 port map( G => n12154, D => N2311, Q 
                           => NEXT_REGISTERS_30_11_port);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => N97, CK => CLK, Q => n_2012
                           , QN => n1973_port);
   NEXT_REGISTERS_reg_30_10_inst : DLH_X1 port map( G => n12153, D => N2310, Q 
                           => NEXT_REGISTERS_30_10_port);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => N96, CK => CLK, Q => n_2013
                           , QN => n1974_port);
   NEXT_REGISTERS_reg_30_9_inst : DLH_X1 port map( G => n12153, D => N2309, Q 
                           => NEXT_REGISTERS_30_9_port);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => N95, CK => CLK, Q => n_2014,
                           QN => n1975_port);
   NEXT_REGISTERS_reg_30_8_inst : DLH_X1 port map( G => n12153, D => N2308, Q 
                           => NEXT_REGISTERS_30_8_port);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => N94, CK => CLK, Q => n_2015,
                           QN => n1976_port);
   NEXT_REGISTERS_reg_30_7_inst : DLH_X1 port map( G => n12153, D => N2307, Q 
                           => NEXT_REGISTERS_30_7_port);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => N93, CK => CLK, Q => n_2016,
                           QN => n1977_port);
   NEXT_REGISTERS_reg_30_6_inst : DLH_X1 port map( G => n12153, D => N2306, Q 
                           => NEXT_REGISTERS_30_6_port);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => N92, CK => CLK, Q => n_2017,
                           QN => n1978_port);
   NEXT_REGISTERS_reg_30_5_inst : DLH_X1 port map( G => n12153, D => N2305, Q 
                           => NEXT_REGISTERS_30_5_port);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => N91, CK => CLK, Q => n_2018,
                           QN => n1979_port);
   NEXT_REGISTERS_reg_30_4_inst : DLH_X1 port map( G => n12153, D => N2304, Q 
                           => NEXT_REGISTERS_30_4_port);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => N90, CK => CLK, Q => n_2019,
                           QN => n1980_port);
   NEXT_REGISTERS_reg_30_3_inst : DLH_X1 port map( G => n12153, D => N2303, Q 
                           => NEXT_REGISTERS_30_3_port);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => N89, CK => CLK, Q => n_2020,
                           QN => n1981_port);
   NEXT_REGISTERS_reg_30_2_inst : DLH_X1 port map( G => n12153, D => N2302, Q 
                           => NEXT_REGISTERS_30_2_port);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => N88, CK => CLK, Q => n_2021,
                           QN => n1982_port);
   NEXT_REGISTERS_reg_30_1_inst : DLH_X1 port map( G => n12153, D => N2301, Q 
                           => NEXT_REGISTERS_30_1_port);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => N87, CK => CLK, Q => n_2022,
                           QN => n1983_port);
   NEXT_REGISTERS_reg_30_0_inst : DLH_X1 port map( G => n12153, D => N2300, Q 
                           => NEXT_REGISTERS_30_0_port);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => N86, CK => CLK, Q => n_2023,
                           QN => n1984_port);
   NEXT_REGISTERS_reg_31_63_inst : DLH_X1 port map( G => n12167, D => N2298, Q 
                           => NEXT_REGISTERS_31_63_port);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => N85, CK => CLK, Q => n_2024
                           , QN => n1985_port);
   NEXT_REGISTERS_reg_31_62_inst : DLH_X1 port map( G => n12167, D => N2297, Q 
                           => NEXT_REGISTERS_31_62_port);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => N84, CK => CLK, Q => n_2025
                           , QN => n1986_port);
   NEXT_REGISTERS_reg_31_61_inst : DLH_X1 port map( G => n12167, D => N2296, Q 
                           => NEXT_REGISTERS_31_61_port);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => N83, CK => CLK, Q => n_2026
                           , QN => n1987_port);
   NEXT_REGISTERS_reg_31_60_inst : DLH_X1 port map( G => n12167, D => N2295, Q 
                           => NEXT_REGISTERS_31_60_port);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => N82, CK => CLK, Q => n_2027
                           , QN => n1988_port);
   NEXT_REGISTERS_reg_31_59_inst : DLH_X1 port map( G => n12167, D => N2294, Q 
                           => NEXT_REGISTERS_31_59_port);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => N81, CK => CLK, Q => n_2028
                           , QN => n1989_port);
   NEXT_REGISTERS_reg_31_58_inst : DLH_X1 port map( G => n12167, D => N2293, Q 
                           => NEXT_REGISTERS_31_58_port);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => N80, CK => CLK, Q => n_2029
                           , QN => n1990_port);
   NEXT_REGISTERS_reg_31_57_inst : DLH_X1 port map( G => n12167, D => N2292, Q 
                           => NEXT_REGISTERS_31_57_port);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => N79, CK => CLK, Q => n_2030
                           , QN => n1991_port);
   NEXT_REGISTERS_reg_31_56_inst : DLH_X1 port map( G => n12167, D => N2291, Q 
                           => NEXT_REGISTERS_31_56_port);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => N78, CK => CLK, Q => n_2031
                           , QN => n1992_port);
   NEXT_REGISTERS_reg_31_55_inst : DLH_X1 port map( G => n12167, D => N2290, Q 
                           => NEXT_REGISTERS_31_55_port);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => N77, CK => CLK, Q => n_2032
                           , QN => n1993_port);
   NEXT_REGISTERS_reg_31_54_inst : DLH_X1 port map( G => n12166, D => N2289, Q 
                           => NEXT_REGISTERS_31_54_port);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => N76, CK => CLK, Q => n_2033
                           , QN => n1994_port);
   NEXT_REGISTERS_reg_31_53_inst : DLH_X1 port map( G => n12166, D => N2288, Q 
                           => NEXT_REGISTERS_31_53_port);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => N75, CK => CLK, Q => n_2034
                           , QN => n1995_port);
   NEXT_REGISTERS_reg_31_52_inst : DLH_X1 port map( G => n12166, D => N2287, Q 
                           => NEXT_REGISTERS_31_52_port);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => N74, CK => CLK, Q => n_2035
                           , QN => n1996_port);
   NEXT_REGISTERS_reg_31_51_inst : DLH_X1 port map( G => n12166, D => N2286, Q 
                           => NEXT_REGISTERS_31_51_port);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => N73, CK => CLK, Q => n_2036
                           , QN => n1997_port);
   NEXT_REGISTERS_reg_31_50_inst : DLH_X1 port map( G => n12166, D => N2285, Q 
                           => NEXT_REGISTERS_31_50_port);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => N72, CK => CLK, Q => n_2037
                           , QN => n1998_port);
   NEXT_REGISTERS_reg_31_49_inst : DLH_X1 port map( G => n12166, D => N2284, Q 
                           => NEXT_REGISTERS_31_49_port);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => N71, CK => CLK, Q => n_2038
                           , QN => n1999_port);
   NEXT_REGISTERS_reg_31_48_inst : DLH_X1 port map( G => n12166, D => N2283, Q 
                           => NEXT_REGISTERS_31_48_port);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => N70, CK => CLK, Q => n_2039
                           , QN => n2000_port);
   NEXT_REGISTERS_reg_31_47_inst : DLH_X1 port map( G => n12166, D => N2282, Q 
                           => NEXT_REGISTERS_31_47_port);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => N69, CK => CLK, Q => n_2040
                           , QN => n2001_port);
   NEXT_REGISTERS_reg_31_46_inst : DLH_X1 port map( G => n12166, D => N2281, Q 
                           => NEXT_REGISTERS_31_46_port);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => N68, CK => CLK, Q => n_2041
                           , QN => n2002_port);
   NEXT_REGISTERS_reg_31_45_inst : DLH_X1 port map( G => n12166, D => N2280, Q 
                           => NEXT_REGISTERS_31_45_port);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => N67, CK => CLK, Q => n_2042
                           , QN => n2003_port);
   NEXT_REGISTERS_reg_31_44_inst : DLH_X1 port map( G => n12166, D => N2279, Q 
                           => NEXT_REGISTERS_31_44_port);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => N66, CK => CLK, Q => n_2043
                           , QN => n2004_port);
   NEXT_REGISTERS_reg_31_43_inst : DLH_X1 port map( G => n12165, D => N2278, Q 
                           => NEXT_REGISTERS_31_43_port);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => N65, CK => CLK, Q => n_2044
                           , QN => n2005_port);
   NEXT_REGISTERS_reg_31_42_inst : DLH_X1 port map( G => n12165, D => N2277, Q 
                           => NEXT_REGISTERS_31_42_port);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => N64, CK => CLK, Q => n_2045
                           , QN => n2006_port);
   NEXT_REGISTERS_reg_31_41_inst : DLH_X1 port map( G => n12165, D => N2276, Q 
                           => NEXT_REGISTERS_31_41_port);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => N63, CK => CLK, Q => n_2046
                           , QN => n2007_port);
   NEXT_REGISTERS_reg_31_40_inst : DLH_X1 port map( G => n12165, D => N2275, Q 
                           => NEXT_REGISTERS_31_40_port);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => N62, CK => CLK, Q => n_2047
                           , QN => n2008_port);
   NEXT_REGISTERS_reg_31_39_inst : DLH_X1 port map( G => n12165, D => N2274, Q 
                           => NEXT_REGISTERS_31_39_port);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => N61, CK => CLK, Q => n_2048
                           , QN => n2009_port);
   NEXT_REGISTERS_reg_31_38_inst : DLH_X1 port map( G => n12165, D => N2273, Q 
                           => NEXT_REGISTERS_31_38_port);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => N60, CK => CLK, Q => n_2049
                           , QN => n2010_port);
   NEXT_REGISTERS_reg_31_37_inst : DLH_X1 port map( G => n12165, D => N2272, Q 
                           => NEXT_REGISTERS_31_37_port);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => N59, CK => CLK, Q => n_2050
                           , QN => n2011_port);
   NEXT_REGISTERS_reg_31_36_inst : DLH_X1 port map( G => n12165, D => N2271, Q 
                           => NEXT_REGISTERS_31_36_port);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => N58, CK => CLK, Q => n_2051
                           , QN => n2012_port);
   NEXT_REGISTERS_reg_31_35_inst : DLH_X1 port map( G => n12165, D => N2270, Q 
                           => NEXT_REGISTERS_31_35_port);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => N57, CK => CLK, Q => n_2052
                           , QN => n2013_port);
   NEXT_REGISTERS_reg_31_34_inst : DLH_X1 port map( G => n12165, D => N2269, Q 
                           => NEXT_REGISTERS_31_34_port);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => N56, CK => CLK, Q => n_2053
                           , QN => n2014_port);
   NEXT_REGISTERS_reg_31_33_inst : DLH_X1 port map( G => n12165, D => N2268, Q 
                           => NEXT_REGISTERS_31_33_port);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => N55, CK => CLK, Q => n_2054
                           , QN => n2015_port);
   NEXT_REGISTERS_reg_31_32_inst : DLH_X1 port map( G => n12164, D => N2267, Q 
                           => NEXT_REGISTERS_31_32_port);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => N54, CK => CLK, Q => n_2055
                           , QN => n2016_port);
   NEXT_REGISTERS_reg_31_31_inst : DLH_X1 port map( G => n12164, D => N2266, Q 
                           => NEXT_REGISTERS_31_31_port);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => N53, CK => CLK, Q => n_2056
                           , QN => n2017_port);
   NEXT_REGISTERS_reg_31_30_inst : DLH_X1 port map( G => n12164, D => N2265, Q 
                           => NEXT_REGISTERS_31_30_port);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => N52, CK => CLK, Q => n_2057
                           , QN => n2018_port);
   NEXT_REGISTERS_reg_31_29_inst : DLH_X1 port map( G => n12164, D => N2264, Q 
                           => NEXT_REGISTERS_31_29_port);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => N51, CK => CLK, Q => n_2058
                           , QN => n2019_port);
   NEXT_REGISTERS_reg_31_28_inst : DLH_X1 port map( G => n12164, D => N2263, Q 
                           => NEXT_REGISTERS_31_28_port);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => N50, CK => CLK, Q => n_2059
                           , QN => n2020_port);
   NEXT_REGISTERS_reg_31_27_inst : DLH_X1 port map( G => n12164, D => N2262, Q 
                           => NEXT_REGISTERS_31_27_port);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => N49, CK => CLK, Q => n_2060
                           , QN => n2021_port);
   NEXT_REGISTERS_reg_31_26_inst : DLH_X1 port map( G => n12164, D => N2261, Q 
                           => NEXT_REGISTERS_31_26_port);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => N48, CK => CLK, Q => n_2061
                           , QN => n2022_port);
   NEXT_REGISTERS_reg_31_25_inst : DLH_X1 port map( G => n12164, D => N2260, Q 
                           => NEXT_REGISTERS_31_25_port);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => N47, CK => CLK, Q => n_2062
                           , QN => n2023_port);
   NEXT_REGISTERS_reg_31_24_inst : DLH_X1 port map( G => n12164, D => N2259, Q 
                           => NEXT_REGISTERS_31_24_port);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => N46, CK => CLK, Q => n_2063
                           , QN => n2024_port);
   NEXT_REGISTERS_reg_31_23_inst : DLH_X1 port map( G => n12164, D => N2258, Q 
                           => NEXT_REGISTERS_31_23_port);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => N45, CK => CLK, Q => n_2064
                           , QN => n2025_port);
   NEXT_REGISTERS_reg_31_22_inst : DLH_X1 port map( G => n12164, D => N2257, Q 
                           => NEXT_REGISTERS_31_22_port);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => N44, CK => CLK, Q => n_2065
                           , QN => n2026_port);
   NEXT_REGISTERS_reg_31_21_inst : DLH_X1 port map( G => n12163, D => N2256, Q 
                           => NEXT_REGISTERS_31_21_port);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => N43, CK => CLK, Q => n_2066
                           , QN => n2027_port);
   NEXT_REGISTERS_reg_31_20_inst : DLH_X1 port map( G => n12163, D => N2255, Q 
                           => NEXT_REGISTERS_31_20_port);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => N42, CK => CLK, Q => n_2067
                           , QN => n2028_port);
   NEXT_REGISTERS_reg_31_19_inst : DLH_X1 port map( G => n12163, D => N2254, Q 
                           => NEXT_REGISTERS_31_19_port);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => N41, CK => CLK, Q => n_2068
                           , QN => n2029_port);
   NEXT_REGISTERS_reg_31_18_inst : DLH_X1 port map( G => n12163, D => N2253, Q 
                           => NEXT_REGISTERS_31_18_port);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => N40, CK => CLK, Q => n_2069
                           , QN => n2030_port);
   NEXT_REGISTERS_reg_31_17_inst : DLH_X1 port map( G => n12163, D => N2252, Q 
                           => NEXT_REGISTERS_31_17_port);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => N39, CK => CLK, Q => n_2070
                           , QN => n2031_port);
   NEXT_REGISTERS_reg_31_16_inst : DLH_X1 port map( G => n12163, D => N2251, Q 
                           => NEXT_REGISTERS_31_16_port);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => N38, CK => CLK, Q => n_2071
                           , QN => n2032_port);
   NEXT_REGISTERS_reg_31_15_inst : DLH_X1 port map( G => n12163, D => N2250, Q 
                           => NEXT_REGISTERS_31_15_port);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => N37, CK => CLK, Q => n_2072
                           , QN => n2033_port);
   NEXT_REGISTERS_reg_31_14_inst : DLH_X1 port map( G => n12163, D => N2249, Q 
                           => NEXT_REGISTERS_31_14_port);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => N36, CK => CLK, Q => n_2073
                           , QN => n2034_port);
   NEXT_REGISTERS_reg_31_13_inst : DLH_X1 port map( G => n12163, D => N2248, Q 
                           => NEXT_REGISTERS_31_13_port);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => N35, CK => CLK, Q => n_2074
                           , QN => n2035_port);
   NEXT_REGISTERS_reg_31_12_inst : DLH_X1 port map( G => n12163, D => N2247, Q 
                           => NEXT_REGISTERS_31_12_port);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => N34, CK => CLK, Q => n_2075
                           , QN => n2036_port);
   NEXT_REGISTERS_reg_31_11_inst : DLH_X1 port map( G => n12163, D => N2246, Q 
                           => NEXT_REGISTERS_31_11_port);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => N33, CK => CLK, Q => n_2076
                           , QN => n2037_port);
   NEXT_REGISTERS_reg_31_10_inst : DLH_X1 port map( G => n12162, D => N2245, Q 
                           => NEXT_REGISTERS_31_10_port);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => N32, CK => CLK, Q => n_2077
                           , QN => n2038_port);
   NEXT_REGISTERS_reg_31_9_inst : DLH_X1 port map( G => n12162, D => N2244, Q 
                           => NEXT_REGISTERS_31_9_port);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => N31, CK => CLK, Q => n_2078,
                           QN => n2039_port);
   NEXT_REGISTERS_reg_31_8_inst : DLH_X1 port map( G => n12162, D => N2243, Q 
                           => NEXT_REGISTERS_31_8_port);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => N30, CK => CLK, Q => n_2079,
                           QN => n2040_port);
   NEXT_REGISTERS_reg_31_7_inst : DLH_X1 port map( G => n12162, D => N2242, Q 
                           => NEXT_REGISTERS_31_7_port);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => N29, CK => CLK, Q => n_2080,
                           QN => n2041_port);
   NEXT_REGISTERS_reg_31_6_inst : DLH_X1 port map( G => n12162, D => N2241, Q 
                           => NEXT_REGISTERS_31_6_port);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => N28, CK => CLK, Q => n_2081,
                           QN => n2042_port);
   NEXT_REGISTERS_reg_31_5_inst : DLH_X1 port map( G => n12162, D => N2240, Q 
                           => NEXT_REGISTERS_31_5_port);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => N27, CK => CLK, Q => n_2082,
                           QN => n2043_port);
   NEXT_REGISTERS_reg_31_4_inst : DLH_X1 port map( G => n12162, D => N2239, Q 
                           => NEXT_REGISTERS_31_4_port);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => N26, CK => CLK, Q => n_2083,
                           QN => n2044_port);
   NEXT_REGISTERS_reg_31_3_inst : DLH_X1 port map( G => n12162, D => N2238, Q 
                           => NEXT_REGISTERS_31_3_port);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => N25, CK => CLK, Q => n_2084,
                           QN => n2045_port);
   NEXT_REGISTERS_reg_31_2_inst : DLH_X1 port map( G => n12162, D => N2237, Q 
                           => NEXT_REGISTERS_31_2_port);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => N24, CK => CLK, Q => n_2085,
                           QN => n2046_port);
   NEXT_REGISTERS_reg_31_1_inst : DLH_X1 port map( G => n12162, D => N2236, Q 
                           => NEXT_REGISTERS_31_1_port);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => N23, CK => CLK, Q => n_2086,
                           QN => n2047_port);
   NEXT_REGISTERS_reg_31_0_inst : DLH_X1 port map( G => n12162, D => N2235, Q 
                           => NEXT_REGISTERS_31_0_port);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => N22, CK => CLK, Q => n_2087,
                           QN => n2048_port);
   U11759 : NAND3_X1 port map( A1 => n6230, A2 => n6229, A3 => n6231, ZN => 
                           n7276);
   U11760 : NAND3_X1 port map( A1 => n6230, A2 => n6229, A3 => ADD_WR(0), ZN =>
                           n7277);
   U11761 : NAND3_X1 port map( A1 => n6231, A2 => n6229, A3 => ADD_WR(1), ZN =>
                           n7278);
   U11762 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n6229, A3 => ADD_WR(1), 
                           ZN => n7279);
   U11763 : NAND3_X1 port map( A1 => n6231, A2 => n6230, A3 => ADD_WR(2), ZN =>
                           n7280);
   U11764 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n6230, A3 => ADD_WR(2), 
                           ZN => n7281);
   U11765 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n6231, A3 => ADD_WR(2), 
                           ZN => n7282);
   U11766 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => 
                           ADD_WR(2), ZN => n7283);
   U11767 : NAND3_X1 port map( A1 => n7287, A2 => n7288, A3 => n7289, ZN => 
                           N2199);
   U11768 : NAND3_X1 port map( A1 => n7327, A2 => n7328, A3 => n7329, ZN => 
                           N2198);
   U11769 : NAND3_X1 port map( A1 => n7345, A2 => n7346, A3 => n7347, ZN => 
                           N2197);
   U11770 : NAND3_X1 port map( A1 => n7363, A2 => n7364, A3 => n7365, ZN => 
                           N2196);
   U11771 : NAND3_X1 port map( A1 => n7381, A2 => n7382, A3 => n7383, ZN => 
                           N2195);
   U11772 : NAND3_X1 port map( A1 => n7399, A2 => n7400, A3 => n7401, ZN => 
                           N2194);
   U11773 : NAND3_X1 port map( A1 => n7417, A2 => n7418, A3 => n7419, ZN => 
                           N2193);
   U11774 : NAND3_X1 port map( A1 => n7435, A2 => n7436, A3 => n7437, ZN => 
                           N2192);
   U11775 : NAND3_X1 port map( A1 => n7453, A2 => n7454, A3 => n7455, ZN => 
                           N2191);
   U11776 : NAND3_X1 port map( A1 => n7471, A2 => n7472, A3 => n7473, ZN => 
                           N2190);
   U11777 : NAND3_X1 port map( A1 => n7489, A2 => n7490, A3 => n7491, ZN => 
                           N2189);
   U11778 : NAND3_X1 port map( A1 => n7507, A2 => n7508, A3 => n7509, ZN => 
                           N2188);
   U11779 : NAND3_X1 port map( A1 => n7525, A2 => n7526, A3 => n7527, ZN => 
                           N2187);
   U11780 : NAND3_X1 port map( A1 => n7543, A2 => n7544, A3 => n7545, ZN => 
                           N2186);
   U11781 : NAND3_X1 port map( A1 => n7561, A2 => n7562, A3 => n7563, ZN => 
                           N2185);
   U11782 : NAND3_X1 port map( A1 => n7579, A2 => n7580, A3 => n7581, ZN => 
                           N2184);
   U11783 : NAND3_X1 port map( A1 => n7597, A2 => n7598, A3 => n7599, ZN => 
                           N2183);
   U11784 : NAND3_X1 port map( A1 => n7615, A2 => n7616, A3 => n7617, ZN => 
                           N2182);
   U11785 : NAND3_X1 port map( A1 => n7633, A2 => n7634, A3 => n7635, ZN => 
                           N2181);
   U11786 : NAND3_X1 port map( A1 => n7651, A2 => n7652, A3 => n7653, ZN => 
                           N2180);
   U11787 : NAND3_X1 port map( A1 => n7669, A2 => n7670, A3 => n7671, ZN => 
                           N2179);
   U11788 : NAND3_X1 port map( A1 => n7687, A2 => n7688, A3 => n7689, ZN => 
                           N2178);
   U11789 : NAND3_X1 port map( A1 => n7705, A2 => n7706, A3 => n7707, ZN => 
                           N2177);
   U11790 : NAND3_X1 port map( A1 => n7723, A2 => n7724, A3 => n7725, ZN => 
                           N2176);
   U11791 : NAND3_X1 port map( A1 => n7741, A2 => n7742, A3 => n7743, ZN => 
                           N2175);
   U11792 : NAND3_X1 port map( A1 => n7759, A2 => n7760, A3 => n7761, ZN => 
                           N2174);
   U11793 : NAND3_X1 port map( A1 => n7777, A2 => n7778, A3 => n7779, ZN => 
                           N2173);
   U11794 : NAND3_X1 port map( A1 => n7795, A2 => n7796, A3 => n7797, ZN => 
                           N2172);
   U11795 : NAND3_X1 port map( A1 => n7813, A2 => n7814, A3 => n7815, ZN => 
                           N2171);
   U11796 : NAND3_X1 port map( A1 => n7831, A2 => n7832, A3 => n7833, ZN => 
                           N2170);
   U11797 : NAND3_X1 port map( A1 => n7849, A2 => n7850, A3 => n7851, ZN => 
                           N2169);
   U11798 : NAND3_X1 port map( A1 => n7867, A2 => n7868, A3 => n7869, ZN => 
                           N2168);
   U11799 : NAND3_X1 port map( A1 => n7885, A2 => n7886, A3 => n7887, ZN => 
                           N2167);
   U11800 : NAND3_X1 port map( A1 => n7903, A2 => n7904, A3 => n7905, ZN => 
                           N2166);
   U11801 : NAND3_X1 port map( A1 => n7921, A2 => n7922, A3 => n7923, ZN => 
                           N2165);
   U11802 : NAND3_X1 port map( A1 => n7939, A2 => n7940, A3 => n7941, ZN => 
                           N2164);
   U11803 : NAND3_X1 port map( A1 => n7957, A2 => n7958, A3 => n7959, ZN => 
                           N2163);
   U11804 : NAND3_X1 port map( A1 => n7975, A2 => n7976, A3 => n7977, ZN => 
                           N2162);
   U11805 : NAND3_X1 port map( A1 => n7993, A2 => n7994, A3 => n7995, ZN => 
                           N2161);
   U11806 : NAND3_X1 port map( A1 => n8011, A2 => n8012, A3 => n8013, ZN => 
                           N2160);
   U11807 : NAND3_X1 port map( A1 => n8029, A2 => n8030, A3 => n8031, ZN => 
                           N2159);
   U11808 : NAND3_X1 port map( A1 => n8047, A2 => n8048, A3 => n8049, ZN => 
                           N2158);
   U11809 : NAND3_X1 port map( A1 => n8065, A2 => n8066, A3 => n8067, ZN => 
                           N2157);
   U11810 : NAND3_X1 port map( A1 => n8083, A2 => n8084, A3 => n8085, ZN => 
                           N2156);
   U11811 : NAND3_X1 port map( A1 => n8101, A2 => n8102, A3 => n8103, ZN => 
                           N2155);
   U11812 : NAND3_X1 port map( A1 => n8119, A2 => n8120, A3 => n8121, ZN => 
                           N2154);
   U11813 : NAND3_X1 port map( A1 => n8137, A2 => n8138, A3 => n8139, ZN => 
                           N2153);
   U11814 : NAND3_X1 port map( A1 => n8155, A2 => n8156, A3 => n8157, ZN => 
                           N2152);
   U11815 : NAND3_X1 port map( A1 => n8173, A2 => n8174, A3 => n8175, ZN => 
                           N2151);
   U11816 : NAND3_X1 port map( A1 => n8191, A2 => n8192, A3 => n8193, ZN => 
                           N2150);
   U11817 : NAND3_X1 port map( A1 => n8209, A2 => n8210, A3 => n8211, ZN => 
                           N2149);
   U11818 : NAND3_X1 port map( A1 => n8227, A2 => n8228, A3 => n8229, ZN => 
                           N2148);
   U11819 : NAND3_X1 port map( A1 => n8245, A2 => n8246, A3 => n8247, ZN => 
                           N2147);
   U11820 : NAND3_X1 port map( A1 => n8263, A2 => n8264, A3 => n8265, ZN => 
                           N2146);
   U11821 : NAND3_X1 port map( A1 => n8281, A2 => n8282, A3 => n8283, ZN => 
                           N2145);
   U11822 : NAND3_X1 port map( A1 => n8299, A2 => n8300, A3 => n8301, ZN => 
                           N2144);
   U11823 : NAND3_X1 port map( A1 => n8317, A2 => n8318, A3 => n8319, ZN => 
                           N2143);
   U11824 : NAND3_X1 port map( A1 => n8335, A2 => n8336, A3 => n8337, ZN => 
                           N2142);
   U11825 : NAND3_X1 port map( A1 => n8353, A2 => n8354, A3 => n8355, ZN => 
                           N2141);
   U11826 : NAND3_X1 port map( A1 => n8371, A2 => n8372, A3 => n8373, ZN => 
                           N2140);
   U11827 : NAND3_X1 port map( A1 => n8389, A2 => n8390, A3 => n8391, ZN => 
                           N2139);
   U11828 : NAND3_X1 port map( A1 => n8407, A2 => n8408, A3 => n8409, ZN => 
                           N2138);
   U11829 : NAND3_X1 port map( A1 => n8425, A2 => n8426, A3 => n8427, ZN => 
                           N2137);
   U11830 : NAND3_X1 port map( A1 => n8443, A2 => n8444, A3 => n8445, ZN => 
                           N2136);
   U11831 : NAND3_X1 port map( A1 => n8467, A2 => n8468, A3 => n8469, ZN => 
                           N2134);
   U11832 : NAND3_X1 port map( A1 => n8507, A2 => n8508, A3 => n8509, ZN => 
                           N2133);
   U11833 : NAND3_X1 port map( A1 => n8525, A2 => n8526, A3 => n8527, ZN => 
                           N2132);
   U11834 : NAND3_X1 port map( A1 => n8543, A2 => n8544, A3 => n8545, ZN => 
                           N2131);
   U11835 : NAND3_X1 port map( A1 => n8561, A2 => n8562, A3 => n8563, ZN => 
                           N2130);
   U11836 : NAND3_X1 port map( A1 => n8579, A2 => n8580, A3 => n8581, ZN => 
                           N2129);
   U11837 : NAND3_X1 port map( A1 => n8597, A2 => n8598, A3 => n8599, ZN => 
                           N2128);
   U11838 : NAND3_X1 port map( A1 => n8615, A2 => n8616, A3 => n8617, ZN => 
                           N2127);
   U11839 : NAND3_X1 port map( A1 => n8633, A2 => n8634, A3 => n8635, ZN => 
                           N2126);
   U11840 : NAND3_X1 port map( A1 => n8651, A2 => n8652, A3 => n8653, ZN => 
                           N2125);
   U11841 : NAND3_X1 port map( A1 => n8669, A2 => n8670, A3 => n8671, ZN => 
                           N2124);
   U11842 : NAND3_X1 port map( A1 => n8687, A2 => n8688, A3 => n8689, ZN => 
                           N2123);
   U11843 : NAND3_X1 port map( A1 => n8705, A2 => n8706, A3 => n8707, ZN => 
                           N2122);
   U11844 : NAND3_X1 port map( A1 => n8723, A2 => n8724, A3 => n8725, ZN => 
                           N2121);
   U11845 : NAND3_X1 port map( A1 => n8741, A2 => n8742, A3 => n8743, ZN => 
                           N2120);
   U11846 : NAND3_X1 port map( A1 => n8759, A2 => n8760, A3 => n8761, ZN => 
                           N2119);
   U11847 : NAND3_X1 port map( A1 => n8777, A2 => n8778, A3 => n8779, ZN => 
                           N2118);
   U11848 : NAND3_X1 port map( A1 => n8795, A2 => n8796, A3 => n8797, ZN => 
                           N2117);
   U11849 : NAND3_X1 port map( A1 => n8813, A2 => n8814, A3 => n8815, ZN => 
                           N2116);
   U11850 : NAND3_X1 port map( A1 => n8831, A2 => n8832, A3 => n8833, ZN => 
                           N2115);
   U11851 : NAND3_X1 port map( A1 => n8849, A2 => n8850, A3 => n8851, ZN => 
                           N2114);
   U11852 : NAND3_X1 port map( A1 => n8867, A2 => n8868, A3 => n8869, ZN => 
                           N2113);
   U11853 : NAND3_X1 port map( A1 => n8885, A2 => n8886, A3 => n8887, ZN => 
                           N2112);
   U11854 : NAND3_X1 port map( A1 => n8903, A2 => n8904, A3 => n8905, ZN => 
                           N2111);
   U11855 : NAND3_X1 port map( A1 => n8921, A2 => n8922, A3 => n8923, ZN => 
                           N2110);
   U11856 : NAND3_X1 port map( A1 => n8939, A2 => n8940, A3 => n8941, ZN => 
                           N2109);
   U11857 : NAND3_X1 port map( A1 => n8957, A2 => n8958, A3 => n8959, ZN => 
                           N2108);
   U11858 : NAND3_X1 port map( A1 => n8975, A2 => n8976, A3 => n8977, ZN => 
                           N2107);
   U11859 : NAND3_X1 port map( A1 => n8993, A2 => n8994, A3 => n8995, ZN => 
                           N2106);
   U11860 : NAND3_X1 port map( A1 => n9011, A2 => n9012, A3 => n9013, ZN => 
                           N2105);
   U11861 : NAND3_X1 port map( A1 => n9029, A2 => n9030, A3 => n9031, ZN => 
                           N2104);
   U11862 : NAND3_X1 port map( A1 => n9047, A2 => n9048, A3 => n9049, ZN => 
                           N2103);
   U11863 : NAND3_X1 port map( A1 => n9065, A2 => n9066, A3 => n9067, ZN => 
                           N2102);
   U11864 : NAND3_X1 port map( A1 => n9083, A2 => n9084, A3 => n9085, ZN => 
                           N2101);
   U11865 : NAND3_X1 port map( A1 => n9101, A2 => n9102, A3 => n9103, ZN => 
                           N2100);
   U11866 : NAND3_X1 port map( A1 => n9119, A2 => n9120, A3 => n9121, ZN => 
                           N2099);
   U11867 : NAND3_X1 port map( A1 => n9137, A2 => n9138, A3 => n9139, ZN => 
                           N2098);
   U11868 : NAND3_X1 port map( A1 => n9155, A2 => n9156, A3 => n9157, ZN => 
                           N2097);
   U11869 : NAND3_X1 port map( A1 => n9173, A2 => n9174, A3 => n9175, ZN => 
                           N2096);
   U11870 : NAND3_X1 port map( A1 => n9191, A2 => n9192, A3 => n9193, ZN => 
                           N2095);
   U11871 : NAND3_X1 port map( A1 => n9209, A2 => n9210, A3 => n9211, ZN => 
                           N2094);
   U11872 : NAND3_X1 port map( A1 => n9227, A2 => n9228, A3 => n9229, ZN => 
                           N2093);
   U11873 : NAND3_X1 port map( A1 => n9245, A2 => n9246, A3 => n9247, ZN => 
                           N2092);
   U11874 : NAND3_X1 port map( A1 => n9263, A2 => n9264, A3 => n9265, ZN => 
                           N2091);
   U11875 : NAND3_X1 port map( A1 => n9281, A2 => n9282, A3 => n9283, ZN => 
                           N2090);
   U11876 : NAND3_X1 port map( A1 => n9299, A2 => n9300, A3 => n9301, ZN => 
                           N2089);
   U11877 : NAND3_X1 port map( A1 => n9317, A2 => n9318, A3 => n9319, ZN => 
                           N2088);
   U11878 : NAND3_X1 port map( A1 => n9335, A2 => n9336, A3 => n9337, ZN => 
                           N2087);
   U11879 : NAND3_X1 port map( A1 => n9353, A2 => n9354, A3 => n9355, ZN => 
                           N2086);
   U11880 : NAND3_X1 port map( A1 => n9371, A2 => n9372, A3 => n9373, ZN => 
                           N2085);
   U11881 : NAND3_X1 port map( A1 => n9389, A2 => n9390, A3 => n9391, ZN => 
                           N2084);
   U11882 : NAND3_X1 port map( A1 => n9407, A2 => n9408, A3 => n9409, ZN => 
                           N2083);
   U11883 : NAND3_X1 port map( A1 => n9425, A2 => n9426, A3 => n9427, ZN => 
                           N2082);
   U11884 : NAND3_X1 port map( A1 => n9443, A2 => n9444, A3 => n9445, ZN => 
                           N2081);
   U11885 : NAND3_X1 port map( A1 => n9461, A2 => n9462, A3 => n9463, ZN => 
                           N2080);
   U11886 : NAND3_X1 port map( A1 => n9479, A2 => n9480, A3 => n9481, ZN => 
                           N2079);
   U11887 : NAND3_X1 port map( A1 => n9497, A2 => n9498, A3 => n9499, ZN => 
                           N2078);
   U11888 : NAND3_X1 port map( A1 => n9515, A2 => n9516, A3 => n9517, ZN => 
                           N2077);
   U11889 : NAND3_X1 port map( A1 => n9533, A2 => n9534, A3 => n9535, ZN => 
                           N2076);
   U11890 : NAND3_X1 port map( A1 => n9551, A2 => n9552, A3 => n9553, ZN => 
                           N2075);
   U11891 : NAND3_X1 port map( A1 => n9569, A2 => n9570, A3 => n9571, ZN => 
                           N2074);
   U11892 : NAND3_X1 port map( A1 => n9587, A2 => n9588, A3 => n9589, ZN => 
                           N2073);
   U11893 : NAND3_X1 port map( A1 => n9605, A2 => n9606, A3 => n9607, ZN => 
                           N2072);
   U11894 : NAND3_X1 port map( A1 => n9623, A2 => n9624, A3 => n9625, ZN => 
                           N2071);
   U11895 : AND2_X1 port map( A1 => n8462, A2 => n11039, ZN => n10607);
   U11896 : AND2_X1 port map( A1 => n9642, A2 => n10814, ZN => n10608);
   U11897 : AND2_X1 port map( A1 => n8462, A2 => n11057, ZN => n10609);
   U11898 : AND2_X1 port map( A1 => n8462, A2 => n8461, ZN => n10610);
   U11899 : AND2_X1 port map( A1 => n8462, A2 => n8460, ZN => n10611);
   U11900 : AND2_X1 port map( A1 => n9642, A2 => n10832, ZN => n10612);
   U11901 : AND2_X1 port map( A1 => n9642, A2 => n9641, ZN => n10613);
   U11902 : AND2_X1 port map( A1 => n9642, A2 => n9640, ZN => n10614);
   U11903 : AND2_X1 port map( A1 => n11021, A2 => n8465, ZN => n10615);
   U11904 : AND2_X1 port map( A1 => n10796, A2 => n9645, ZN => n10616);
   U11905 : AND2_X1 port map( A1 => n8458, A2 => n8465, ZN => n10617);
   U11906 : AND2_X1 port map( A1 => n8460, A2 => n8465, ZN => n10618);
   U11907 : AND2_X1 port map( A1 => n9638, A2 => n9645, ZN => n10619);
   U11908 : AND2_X1 port map( A1 => n9640, A2 => n9645, ZN => n10620);
   U11909 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n10621);
   U11910 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n10622);
   U11911 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n10623);
   U11912 : BUF_X1 port map( A => n10609, Z => n10932);
   U11913 : BUF_X1 port map( A => n10609, Z => n10933);
   U11914 : BUF_X1 port map( A => n10612, Z => n10707);
   U11915 : BUF_X1 port map( A => n10612, Z => n10708);
   U11916 : BUF_X1 port map( A => n10607, Z => n10873);
   U11917 : BUF_X1 port map( A => n10607, Z => n10874);
   U11918 : BUF_X1 port map( A => n10608, Z => n10648);
   U11919 : BUF_X1 port map( A => n10608, Z => n10649);
   U11920 : BUF_X1 port map( A => n10950, Z => n10957);
   U11921 : BUF_X1 port map( A => n10977, Z => n10984);
   U11922 : BUF_X1 port map( A => n10950, Z => n10958);
   U11923 : BUF_X1 port map( A => n10977, Z => n10985);
   U11924 : BUF_X1 port map( A => n10725, Z => n10732);
   U11925 : BUF_X1 port map( A => n10752, Z => n10759);
   U11926 : BUF_X1 port map( A => n10725, Z => n10733);
   U11927 : BUF_X1 port map( A => n10752, Z => n10760);
   U11928 : BUF_X1 port map( A => n11891, Z => n11889);
   U11929 : BUF_X1 port map( A => n11891, Z => n11890);
   U11930 : BUF_X1 port map( A => n11531, Z => n11544);
   U11931 : BUF_X1 port map( A => n11548, Z => n11561);
   U11932 : BUF_X1 port map( A => n11582, Z => n11595);
   U11933 : BUF_X1 port map( A => n11565, Z => n11578);
   U11934 : BUF_X1 port map( A => n11531, Z => n11545);
   U11935 : BUF_X1 port map( A => n11548, Z => n11562);
   U11936 : BUF_X1 port map( A => n11582, Z => n11596);
   U11937 : BUF_X1 port map( A => n11565, Z => n11579);
   U11938 : BUF_X1 port map( A => n11531, Z => n11546);
   U11939 : BUF_X1 port map( A => n11548, Z => n11563);
   U11940 : BUF_X1 port map( A => n11582, Z => n11597);
   U11941 : BUF_X1 port map( A => n11565, Z => n11580);
   U11942 : BUF_X1 port map( A => n11599, Z => n11612);
   U11943 : BUF_X1 port map( A => n11616, Z => n11629);
   U11944 : BUF_X1 port map( A => n11650, Z => n11663);
   U11945 : BUF_X1 port map( A => n11633, Z => n11646);
   U11946 : BUF_X1 port map( A => n11599, Z => n11613);
   U11947 : BUF_X1 port map( A => n11616, Z => n11630);
   U11948 : BUF_X1 port map( A => n11650, Z => n11664);
   U11949 : BUF_X1 port map( A => n11633, Z => n11647);
   U11950 : BUF_X1 port map( A => n11599, Z => n11614);
   U11951 : BUF_X1 port map( A => n11616, Z => n11631);
   U11952 : BUF_X1 port map( A => n11650, Z => n11665);
   U11953 : BUF_X1 port map( A => n11633, Z => n11648);
   U11954 : BUF_X1 port map( A => n11026, Z => n11024);
   U11955 : BUF_X1 port map( A => n11026, Z => n11023);
   U11956 : BUF_X1 port map( A => n10801, Z => n10799);
   U11957 : BUF_X1 port map( A => n10801, Z => n10798);
   U11958 : BUF_X1 port map( A => n11880, Z => n11878);
   U11959 : BUF_X1 port map( A => n11880, Z => n11879);
   U11960 : BUF_X1 port map( A => n11881, Z => n11874);
   U11961 : BUF_X1 port map( A => n11881, Z => n11875);
   U11962 : BUF_X1 port map( A => n11881, Z => n11876);
   U11963 : BUF_X1 port map( A => n11880, Z => n11877);
   U11964 : BUF_X1 port map( A => n6246, Z => n11531);
   U11965 : BUF_X1 port map( A => n6245, Z => n11548);
   U11966 : BUF_X1 port map( A => n6243, Z => n11582);
   U11967 : BUF_X1 port map( A => n6244, Z => n11565);
   U11968 : BUF_X1 port map( A => n6237, Z => n11599);
   U11969 : BUF_X1 port map( A => n6236, Z => n11616);
   U11970 : BUF_X1 port map( A => n6234, Z => n11650);
   U11971 : BUF_X1 port map( A => n6235, Z => n11633);
   U11972 : BUF_X1 port map( A => n11028, Z => n11026);
   U11973 : BUF_X1 port map( A => n10803, Z => n10801);
   U11974 : BUF_X1 port map( A => n10611, Z => n10948);
   U11975 : BUF_X1 port map( A => n10610, Z => n10940);
   U11976 : BUF_X1 port map( A => n10611, Z => n10949);
   U11977 : BUF_X1 port map( A => n10610, Z => n10941);
   U11978 : BUF_X1 port map( A => n10614, Z => n10723);
   U11979 : BUF_X1 port map( A => n10613, Z => n10715);
   U11980 : BUF_X1 port map( A => n10614, Z => n10724);
   U11981 : BUF_X1 port map( A => n10613, Z => n10716);
   U11982 : BUF_X1 port map( A => n10883, Z => n10890);
   U11983 : BUF_X1 port map( A => n10892, Z => n10899);
   U11984 : BUF_X1 port map( A => n10901, Z => n10908);
   U11985 : BUF_X1 port map( A => n10858, Z => n10865);
   U11986 : BUF_X1 port map( A => n10849, Z => n10856);
   U11987 : BUF_X1 port map( A => n10959, Z => n10966);
   U11988 : BUF_X1 port map( A => n10968, Z => n10975);
   U11989 : BUF_X1 port map( A => n11065, Z => n11072);
   U11990 : BUF_X1 port map( A => n10883, Z => n10891);
   U11991 : BUF_X1 port map( A => n10892, Z => n10900);
   U11992 : BUF_X1 port map( A => n10901, Z => n10909);
   U11993 : BUF_X1 port map( A => n10858, Z => n10866);
   U11994 : BUF_X1 port map( A => n10849, Z => n10857);
   U11995 : BUF_X1 port map( A => n10959, Z => n10967);
   U11996 : BUF_X1 port map( A => n10968, Z => n10976);
   U11997 : BUF_X1 port map( A => n11065, Z => n11073);
   U11998 : BUF_X1 port map( A => n10658, Z => n10665);
   U11999 : BUF_X1 port map( A => n10667, Z => n10674);
   U12000 : BUF_X1 port map( A => n10676, Z => n10683);
   U12001 : BUF_X1 port map( A => n10633, Z => n10640);
   U12002 : BUF_X1 port map( A => n10624, Z => n10631);
   U12003 : BUF_X1 port map( A => n10734, Z => n10741);
   U12004 : BUF_X1 port map( A => n10743, Z => n10750);
   U12005 : BUF_X1 port map( A => n10840, Z => n10847);
   U12006 : BUF_X1 port map( A => n10658, Z => n10666);
   U12007 : BUF_X1 port map( A => n10667, Z => n10675);
   U12008 : BUF_X1 port map( A => n10676, Z => n10684);
   U12009 : BUF_X1 port map( A => n10633, Z => n10641);
   U12010 : BUF_X1 port map( A => n10624, Z => n10632);
   U12011 : BUF_X1 port map( A => n10734, Z => n10742);
   U12012 : BUF_X1 port map( A => n10743, Z => n10751);
   U12013 : BUF_X1 port map( A => n10840, Z => n10848);
   U12014 : BUF_X1 port map( A => n11530, Z => n11524);
   U12015 : BUF_X1 port map( A => n11530, Z => n11525);
   U12016 : BUF_X1 port map( A => n10618, Z => n10924);
   U12017 : BUF_X1 port map( A => n10617, Z => n10916);
   U12018 : BUF_X1 port map( A => n10615, Z => n10881);
   U12019 : BUF_X1 port map( A => n10618, Z => n10925);
   U12020 : BUF_X1 port map( A => n10617, Z => n10917);
   U12021 : BUF_X1 port map( A => n10615, Z => n10882);
   U12022 : BUF_X1 port map( A => n10620, Z => n10699);
   U12023 : BUF_X1 port map( A => n10619, Z => n10691);
   U12024 : BUF_X1 port map( A => n10616, Z => n10656);
   U12025 : BUF_X1 port map( A => n10620, Z => n10700);
   U12026 : BUF_X1 port map( A => n10619, Z => n10692);
   U12027 : BUF_X1 port map( A => n10616, Z => n10657);
   U12028 : BUF_X1 port map( A => n12170, Z => n12169);
   U12029 : BUF_X1 port map( A => n12170, Z => n12168);
   U12030 : BUF_X1 port map( A => n12161, Z => n12160);
   U12031 : BUF_X1 port map( A => n12161, Z => n12159);
   U12032 : BUF_X1 port map( A => n12152, Z => n12150);
   U12033 : BUF_X1 port map( A => n12152, Z => n12151);
   U12034 : BUF_X1 port map( A => n12143, Z => n12141);
   U12035 : BUF_X1 port map( A => n12143, Z => n12142);
   U12036 : BUF_X1 port map( A => n12134, Z => n12132);
   U12037 : BUF_X1 port map( A => n12134, Z => n12133);
   U12038 : BUF_X1 port map( A => n12125, Z => n12123);
   U12039 : BUF_X1 port map( A => n12125, Z => n12124);
   U12040 : BUF_X1 port map( A => n12116, Z => n12114);
   U12041 : BUF_X1 port map( A => n12116, Z => n12115);
   U12042 : BUF_X1 port map( A => n12107, Z => n12105);
   U12043 : BUF_X1 port map( A => n12107, Z => n12106);
   U12044 : BUF_X1 port map( A => n12098, Z => n12096);
   U12045 : BUF_X1 port map( A => n12098, Z => n12097);
   U12046 : BUF_X1 port map( A => n12089, Z => n12087);
   U12047 : BUF_X1 port map( A => n12089, Z => n12088);
   U12048 : BUF_X1 port map( A => n12080, Z => n12078);
   U12049 : BUF_X1 port map( A => n12080, Z => n12079);
   U12050 : BUF_X1 port map( A => n12071, Z => n12069);
   U12051 : BUF_X1 port map( A => n12071, Z => n12070);
   U12052 : BUF_X1 port map( A => n12062, Z => n12060);
   U12053 : BUF_X1 port map( A => n12062, Z => n12061);
   U12054 : BUF_X1 port map( A => n12053, Z => n12051);
   U12055 : BUF_X1 port map( A => n12053, Z => n12052);
   U12056 : BUF_X1 port map( A => n12044, Z => n12042);
   U12057 : BUF_X1 port map( A => n12044, Z => n12043);
   U12058 : BUF_X1 port map( A => n12035, Z => n12033);
   U12059 : BUF_X1 port map( A => n12035, Z => n12034);
   U12060 : BUF_X1 port map( A => n12026, Z => n12024);
   U12061 : BUF_X1 port map( A => n12026, Z => n12025);
   U12062 : BUF_X1 port map( A => n12017, Z => n12015);
   U12063 : BUF_X1 port map( A => n12017, Z => n12016);
   U12064 : BUF_X1 port map( A => n12008, Z => n12006);
   U12065 : BUF_X1 port map( A => n12008, Z => n12007);
   U12066 : BUF_X1 port map( A => n11999, Z => n11997);
   U12067 : BUF_X1 port map( A => n11999, Z => n11998);
   U12068 : BUF_X1 port map( A => n11990, Z => n11988);
   U12069 : BUF_X1 port map( A => n11990, Z => n11989);
   U12070 : BUF_X1 port map( A => n11981, Z => n11979);
   U12071 : BUF_X1 port map( A => n11981, Z => n11980);
   U12072 : BUF_X1 port map( A => n11972, Z => n11970);
   U12073 : BUF_X1 port map( A => n11972, Z => n11971);
   U12074 : BUF_X1 port map( A => n11963, Z => n11961);
   U12075 : BUF_X1 port map( A => n11963, Z => n11962);
   U12076 : BUF_X1 port map( A => n11954, Z => n11952);
   U12077 : BUF_X1 port map( A => n11954, Z => n11953);
   U12078 : BUF_X1 port map( A => n11945, Z => n11943);
   U12079 : BUF_X1 port map( A => n11945, Z => n11944);
   U12080 : BUF_X1 port map( A => n11936, Z => n11934);
   U12081 : BUF_X1 port map( A => n11936, Z => n11935);
   U12082 : BUF_X1 port map( A => n11927, Z => n11925);
   U12083 : BUF_X1 port map( A => n11927, Z => n11926);
   U12084 : BUF_X1 port map( A => n11918, Z => n11916);
   U12085 : BUF_X1 port map( A => n11918, Z => n11917);
   U12086 : BUF_X1 port map( A => n11909, Z => n11907);
   U12087 : BUF_X1 port map( A => n11909, Z => n11908);
   U12088 : BUF_X1 port map( A => n11900, Z => n11898);
   U12089 : BUF_X1 port map( A => n11900, Z => n11899);
   U12090 : BUF_X1 port map( A => n11529, Z => n11527);
   U12091 : BUF_X1 port map( A => n11529, Z => n11528);
   U12092 : BUF_X1 port map( A => n11529, Z => n11526);
   U12093 : BUF_X1 port map( A => n11009, Z => n11007);
   U12094 : BUF_X1 port map( A => n11044, Z => n11042);
   U12095 : BUF_X1 port map( A => n11062, Z => n11060);
   U12096 : BUF_X1 port map( A => n11009, Z => n11006);
   U12097 : BUF_X1 port map( A => n11062, Z => n11059);
   U12098 : BUF_X1 port map( A => n11044, Z => n11041);
   U12099 : BUF_X1 port map( A => n10784, Z => n10782);
   U12100 : BUF_X1 port map( A => n10819, Z => n10817);
   U12101 : BUF_X1 port map( A => n10837, Z => n10835);
   U12102 : BUF_X1 port map( A => n10784, Z => n10781);
   U12103 : BUF_X1 port map( A => n10837, Z => n10834);
   U12104 : BUF_X1 port map( A => n10819, Z => n10816);
   U12105 : BUF_X1 port map( A => n11027, Z => n11022);
   U12106 : BUF_X1 port map( A => n10802, Z => n10797);
   U12107 : BUF_X1 port map( A => n11882, Z => n11873);
   U12108 : BUF_X1 port map( A => n10621, Z => n11529);
   U12109 : BUF_X1 port map( A => n6226, Z => n11881);
   U12110 : BUF_X1 port map( A => n6226, Z => n11880);
   U12111 : BUF_X1 port map( A => n11011, Z => n11009);
   U12112 : BUF_X1 port map( A => n11064, Z => n11062);
   U12113 : BUF_X1 port map( A => n11046, Z => n11044);
   U12114 : BUF_X1 port map( A => n10786, Z => n10784);
   U12115 : BUF_X1 port map( A => n10839, Z => n10837);
   U12116 : BUF_X1 port map( A => n10821, Z => n10819);
   U12117 : BUF_X1 port map( A => n10986, Z => n10993);
   U12118 : BUF_X1 port map( A => n10986, Z => n10994);
   U12119 : BUF_X1 port map( A => n10761, Z => n10768);
   U12120 : BUF_X1 port map( A => n10761, Z => n10769);
   U12121 : BUF_X1 port map( A => n10622, Z => n12178);
   U12122 : BUF_X1 port map( A => n10622, Z => n12177);
   U12123 : BUF_X1 port map( A => n10623, Z => n12186);
   U12124 : BUF_X1 port map( A => n10623, Z => n12185);
   U12125 : BUF_X1 port map( A => n11010, Z => n11005);
   U12126 : BUF_X1 port map( A => n11063, Z => n11058);
   U12127 : BUF_X1 port map( A => n11045, Z => n11040);
   U12128 : BUF_X1 port map( A => n10785, Z => n10780);
   U12129 : BUF_X1 port map( A => n10838, Z => n10833);
   U12130 : BUF_X1 port map( A => n10820, Z => n10815);
   U12131 : BUF_X1 port map( A => n7274, Z => n11074);
   U12132 : BUF_X1 port map( A => n7272, Z => n11082);
   U12133 : BUF_X1 port map( A => n7269, Z => n11094);
   U12134 : BUF_X1 port map( A => n7268, Z => n11098);
   U12135 : BUF_X1 port map( A => n7273, Z => n11078);
   U12136 : BUF_X1 port map( A => n7271, Z => n11086);
   U12137 : BUF_X1 port map( A => n7270, Z => n11090);
   U12138 : BUF_X1 port map( A => n7267, Z => n11102);
   U12139 : BUF_X1 port map( A => n7266, Z => n11106);
   U12140 : BUF_X1 port map( A => n7265, Z => n11110);
   U12141 : BUF_X1 port map( A => n7264, Z => n11114);
   U12142 : BUF_X1 port map( A => n7263, Z => n11118);
   U12143 : BUF_X1 port map( A => n7262, Z => n11122);
   U12144 : BUF_X1 port map( A => n7261, Z => n11126);
   U12145 : BUF_X1 port map( A => n7260, Z => n11130);
   U12146 : BUF_X1 port map( A => n7259, Z => n11134);
   U12147 : BUF_X1 port map( A => n7258, Z => n11138);
   U12148 : BUF_X1 port map( A => n7257, Z => n11142);
   U12149 : BUF_X1 port map( A => n7256, Z => n11146);
   U12150 : BUF_X1 port map( A => n7255, Z => n11150);
   U12151 : BUF_X1 port map( A => n7254, Z => n11154);
   U12152 : BUF_X1 port map( A => n7253, Z => n11158);
   U12153 : BUF_X1 port map( A => n7252, Z => n11162);
   U12154 : BUF_X1 port map( A => n7251, Z => n11166);
   U12155 : BUF_X1 port map( A => n7250, Z => n11170);
   U12156 : BUF_X1 port map( A => n7249, Z => n11174);
   U12157 : BUF_X1 port map( A => n7248, Z => n11178);
   U12158 : BUF_X1 port map( A => n7247, Z => n11182);
   U12159 : BUF_X1 port map( A => n7246, Z => n11186);
   U12160 : BUF_X1 port map( A => n7245, Z => n11190);
   U12161 : BUF_X1 port map( A => n7244, Z => n11194);
   U12162 : BUF_X1 port map( A => n7243, Z => n11198);
   U12163 : BUF_X1 port map( A => n7242, Z => n11202);
   U12164 : BUF_X1 port map( A => n7241, Z => n11206);
   U12165 : BUF_X1 port map( A => n7240, Z => n11210);
   U12166 : BUF_X1 port map( A => n7239, Z => n11214);
   U12167 : BUF_X1 port map( A => n7238, Z => n11218);
   U12168 : BUF_X1 port map( A => n7237, Z => n11222);
   U12169 : BUF_X1 port map( A => n7236, Z => n11226);
   U12170 : BUF_X1 port map( A => n7235, Z => n11230);
   U12171 : BUF_X1 port map( A => n7234, Z => n11234);
   U12172 : BUF_X1 port map( A => n7233, Z => n11238);
   U12173 : BUF_X1 port map( A => n7232, Z => n11242);
   U12174 : BUF_X1 port map( A => n7231, Z => n11246);
   U12175 : BUF_X1 port map( A => n7230, Z => n11250);
   U12176 : BUF_X1 port map( A => n7229, Z => n11254);
   U12177 : BUF_X1 port map( A => n7228, Z => n11258);
   U12178 : BUF_X1 port map( A => n7227, Z => n11262);
   U12179 : BUF_X1 port map( A => n7226, Z => n11266);
   U12180 : BUF_X1 port map( A => n7225, Z => n11270);
   U12181 : BUF_X1 port map( A => n7224, Z => n11274);
   U12182 : BUF_X1 port map( A => n7223, Z => n11278);
   U12183 : BUF_X1 port map( A => n7222, Z => n11282);
   U12184 : BUF_X1 port map( A => n7221, Z => n11286);
   U12185 : BUF_X1 port map( A => n7220, Z => n11290);
   U12186 : BUF_X1 port map( A => n7219, Z => n11294);
   U12187 : BUF_X1 port map( A => n7218, Z => n11298);
   U12188 : BUF_X1 port map( A => n7217, Z => n11302);
   U12189 : BUF_X1 port map( A => n7216, Z => n11306);
   U12190 : BUF_X1 port map( A => n7215, Z => n11310);
   U12191 : BUF_X1 port map( A => n7214, Z => n11314);
   U12192 : BUF_X1 port map( A => n7213, Z => n11318);
   U12193 : BUF_X1 port map( A => n7212, Z => n11322);
   U12194 : BUF_X1 port map( A => n7211, Z => n11326);
   U12195 : BUF_X1 port map( A => n11509, Z => n11506);
   U12196 : BUF_X1 port map( A => n11509, Z => n11507);
   U12197 : BUF_X1 port map( A => n11523, Z => n11334);
   U12198 : BUF_X1 port map( A => n11523, Z => n11333);
   U12199 : BUF_X1 port map( A => n11523, Z => n11331);
   U12200 : BUF_X1 port map( A => n11523, Z => n11330);
   U12201 : BUF_X1 port map( A => n11523, Z => n11332);
   U12202 : BUF_X1 port map( A => n11523, Z => n11335);
   U12203 : BUF_X1 port map( A => n11513, Z => n11452);
   U12204 : BUF_X1 port map( A => n11513, Z => n11451);
   U12205 : BUF_X1 port map( A => n11513, Z => n11450);
   U12206 : BUF_X1 port map( A => n11513, Z => n11449);
   U12207 : BUF_X1 port map( A => n11514, Z => n11447);
   U12208 : BUF_X1 port map( A => n11514, Z => n11446);
   U12209 : BUF_X1 port map( A => n11514, Z => n11445);
   U12210 : BUF_X1 port map( A => n11514, Z => n11444);
   U12211 : BUF_X1 port map( A => n11514, Z => n11443);
   U12212 : BUF_X1 port map( A => n11514, Z => n11448);
   U12213 : BUF_X1 port map( A => n11512, Z => n11463);
   U12214 : BUF_X1 port map( A => n11512, Z => n11462);
   U12215 : BUF_X1 port map( A => n11512, Z => n11461);
   U12216 : BUF_X1 port map( A => n11513, Z => n11460);
   U12217 : BUF_X1 port map( A => n11513, Z => n11459);
   U12218 : BUF_X1 port map( A => n11513, Z => n11457);
   U12219 : BUF_X1 port map( A => n11513, Z => n11456);
   U12220 : BUF_X1 port map( A => n11513, Z => n11455);
   U12221 : BUF_X1 port map( A => n11513, Z => n11454);
   U12222 : BUF_X1 port map( A => n11513, Z => n11453);
   U12223 : BUF_X1 port map( A => n11513, Z => n11458);
   U12224 : BUF_X1 port map( A => n11515, Z => n11431);
   U12225 : BUF_X1 port map( A => n11515, Z => n11430);
   U12226 : BUF_X1 port map( A => n11515, Z => n11429);
   U12227 : BUF_X1 port map( A => n11515, Z => n11428);
   U12228 : BUF_X1 port map( A => n11515, Z => n11427);
   U12229 : BUF_X1 port map( A => n11515, Z => n11425);
   U12230 : BUF_X1 port map( A => n11516, Z => n11424);
   U12231 : BUF_X1 port map( A => n11516, Z => n11423);
   U12232 : BUF_X1 port map( A => n11516, Z => n11422);
   U12233 : BUF_X1 port map( A => n11515, Z => n11426);
   U12234 : BUF_X1 port map( A => n11514, Z => n11441);
   U12235 : BUF_X1 port map( A => n11514, Z => n11440);
   U12236 : BUF_X1 port map( A => n11514, Z => n11439);
   U12237 : BUF_X1 port map( A => n11514, Z => n11438);
   U12238 : BUF_X1 port map( A => n11515, Z => n11436);
   U12239 : BUF_X1 port map( A => n11515, Z => n11435);
   U12240 : BUF_X1 port map( A => n11515, Z => n11434);
   U12241 : BUF_X1 port map( A => n11515, Z => n11433);
   U12242 : BUF_X1 port map( A => n11515, Z => n11432);
   U12243 : BUF_X1 port map( A => n11514, Z => n11437);
   U12244 : BUF_X1 port map( A => n11514, Z => n11442);
   U12245 : BUF_X1 port map( A => n11510, Z => n11495);
   U12246 : BUF_X1 port map( A => n11510, Z => n11494);
   U12247 : BUF_X1 port map( A => n11510, Z => n11493);
   U12248 : BUF_X1 port map( A => n11510, Z => n11492);
   U12249 : BUF_X1 port map( A => n11510, Z => n11490);
   U12250 : BUF_X1 port map( A => n11510, Z => n11489);
   U12251 : BUF_X1 port map( A => n11510, Z => n11488);
   U12252 : BUF_X1 port map( A => n11510, Z => n11487);
   U12253 : BUF_X1 port map( A => n11510, Z => n11486);
   U12254 : BUF_X1 port map( A => n11509, Z => n11505);
   U12255 : BUF_X1 port map( A => n11509, Z => n11504);
   U12256 : BUF_X1 port map( A => n11509, Z => n11503);
   U12257 : BUF_X1 port map( A => n11509, Z => n11502);
   U12258 : BUF_X1 port map( A => n11509, Z => n11500);
   U12259 : BUF_X1 port map( A => n11509, Z => n11499);
   U12260 : BUF_X1 port map( A => n11509, Z => n11498);
   U12261 : BUF_X1 port map( A => n11509, Z => n11497);
   U12262 : BUF_X1 port map( A => n11510, Z => n11496);
   U12263 : BUF_X1 port map( A => n11509, Z => n11501);
   U12264 : BUF_X1 port map( A => n11511, Z => n11474);
   U12265 : BUF_X1 port map( A => n11511, Z => n11473);
   U12266 : BUF_X1 port map( A => n11512, Z => n11472);
   U12267 : BUF_X1 port map( A => n11512, Z => n11471);
   U12268 : BUF_X1 port map( A => n11512, Z => n11470);
   U12269 : BUF_X1 port map( A => n11512, Z => n11468);
   U12270 : BUF_X1 port map( A => n11512, Z => n11467);
   U12271 : BUF_X1 port map( A => n11512, Z => n11466);
   U12272 : BUF_X1 port map( A => n11512, Z => n11465);
   U12273 : BUF_X1 port map( A => n11512, Z => n11464);
   U12274 : BUF_X1 port map( A => n11512, Z => n11469);
   U12275 : BUF_X1 port map( A => n11510, Z => n11485);
   U12276 : BUF_X1 port map( A => n11511, Z => n11484);
   U12277 : BUF_X1 port map( A => n11511, Z => n11483);
   U12278 : BUF_X1 port map( A => n11511, Z => n11482);
   U12279 : BUF_X1 port map( A => n11511, Z => n11481);
   U12280 : BUF_X1 port map( A => n11511, Z => n11479);
   U12281 : BUF_X1 port map( A => n11511, Z => n11478);
   U12282 : BUF_X1 port map( A => n11511, Z => n11477);
   U12283 : BUF_X1 port map( A => n11511, Z => n11476);
   U12284 : BUF_X1 port map( A => n11511, Z => n11475);
   U12285 : BUF_X1 port map( A => n11511, Z => n11480);
   U12286 : BUF_X1 port map( A => n11510, Z => n11491);
   U12287 : BUF_X1 port map( A => n11520, Z => n11366);
   U12288 : BUF_X1 port map( A => n11520, Z => n11365);
   U12289 : BUF_X1 port map( A => n11521, Z => n11364);
   U12290 : BUF_X1 port map( A => n11521, Z => n11363);
   U12291 : BUF_X1 port map( A => n11521, Z => n11361);
   U12292 : BUF_X1 port map( A => n11521, Z => n11360);
   U12293 : BUF_X1 port map( A => n11521, Z => n11359);
   U12294 : BUF_X1 port map( A => n11521, Z => n11358);
   U12295 : BUF_X1 port map( A => n11521, Z => n11357);
   U12296 : BUF_X1 port map( A => n11521, Z => n11362);
   U12297 : BUF_X1 port map( A => n11519, Z => n11377);
   U12298 : BUF_X1 port map( A => n11520, Z => n11376);
   U12299 : BUF_X1 port map( A => n11520, Z => n11375);
   U12300 : BUF_X1 port map( A => n11520, Z => n11374);
   U12301 : BUF_X1 port map( A => n11520, Z => n11373);
   U12302 : BUF_X1 port map( A => n11520, Z => n11371);
   U12303 : BUF_X1 port map( A => n11520, Z => n11370);
   U12304 : BUF_X1 port map( A => n11520, Z => n11369);
   U12305 : BUF_X1 port map( A => n11520, Z => n11368);
   U12306 : BUF_X1 port map( A => n11520, Z => n11367);
   U12307 : BUF_X1 port map( A => n11520, Z => n11372);
   U12308 : BUF_X1 port map( A => n11522, Z => n11345);
   U12309 : BUF_X1 port map( A => n11522, Z => n11344);
   U12310 : BUF_X1 port map( A => n11522, Z => n11343);
   U12311 : BUF_X1 port map( A => n11522, Z => n11342);
   U12312 : BUF_X1 port map( A => n11522, Z => n11341);
   U12313 : BUF_X1 port map( A => n11523, Z => n11336);
   U12314 : BUF_X1 port map( A => n11523, Z => n11337);
   U12315 : BUF_X1 port map( A => n11523, Z => n11338);
   U12316 : BUF_X1 port map( A => n11523, Z => n11339);
   U12317 : BUF_X1 port map( A => n11521, Z => n11355);
   U12318 : BUF_X1 port map( A => n11521, Z => n11354);
   U12319 : BUF_X1 port map( A => n11521, Z => n11353);
   U12320 : BUF_X1 port map( A => n11522, Z => n11352);
   U12321 : BUF_X1 port map( A => n11522, Z => n11350);
   U12322 : BUF_X1 port map( A => n11522, Z => n11349);
   U12323 : BUF_X1 port map( A => n11522, Z => n11348);
   U12324 : BUF_X1 port map( A => n11522, Z => n11347);
   U12325 : BUF_X1 port map( A => n11522, Z => n11346);
   U12326 : BUF_X1 port map( A => n11522, Z => n11351);
   U12327 : BUF_X1 port map( A => n11521, Z => n11356);
   U12328 : BUF_X1 port map( A => n11517, Z => n11409);
   U12329 : BUF_X1 port map( A => n11517, Z => n11408);
   U12330 : BUF_X1 port map( A => n11517, Z => n11407);
   U12331 : BUF_X1 port map( A => n11517, Z => n11406);
   U12332 : BUF_X1 port map( A => n11517, Z => n11404);
   U12333 : BUF_X1 port map( A => n11517, Z => n11403);
   U12334 : BUF_X1 port map( A => n11517, Z => n11402);
   U12335 : BUF_X1 port map( A => n11517, Z => n11401);
   U12336 : BUF_X1 port map( A => n11518, Z => n11400);
   U12337 : BUF_X1 port map( A => n11517, Z => n11405);
   U12338 : BUF_X1 port map( A => n11516, Z => n11420);
   U12339 : BUF_X1 port map( A => n11516, Z => n11419);
   U12340 : BUF_X1 port map( A => n11516, Z => n11418);
   U12341 : BUF_X1 port map( A => n11516, Z => n11417);
   U12342 : BUF_X1 port map( A => n11516, Z => n11416);
   U12343 : BUF_X1 port map( A => n11516, Z => n11414);
   U12344 : BUF_X1 port map( A => n11516, Z => n11413);
   U12345 : BUF_X1 port map( A => n11517, Z => n11412);
   U12346 : BUF_X1 port map( A => n11517, Z => n11411);
   U12347 : BUF_X1 port map( A => n11517, Z => n11410);
   U12348 : BUF_X1 port map( A => n11516, Z => n11415);
   U12349 : BUF_X1 port map( A => n11519, Z => n11388);
   U12350 : BUF_X1 port map( A => n11519, Z => n11387);
   U12351 : BUF_X1 port map( A => n11519, Z => n11386);
   U12352 : BUF_X1 port map( A => n11519, Z => n11385);
   U12353 : BUF_X1 port map( A => n11519, Z => n11384);
   U12354 : BUF_X1 port map( A => n11519, Z => n11382);
   U12355 : BUF_X1 port map( A => n11519, Z => n11381);
   U12356 : BUF_X1 port map( A => n11519, Z => n11380);
   U12357 : BUF_X1 port map( A => n11519, Z => n11379);
   U12358 : BUF_X1 port map( A => n11519, Z => n11378);
   U12359 : BUF_X1 port map( A => n11519, Z => n11383);
   U12360 : BUF_X1 port map( A => n11518, Z => n11398);
   U12361 : BUF_X1 port map( A => n11518, Z => n11397);
   U12362 : BUF_X1 port map( A => n11518, Z => n11396);
   U12363 : BUF_X1 port map( A => n11518, Z => n11395);
   U12364 : BUF_X1 port map( A => n11518, Z => n11393);
   U12365 : BUF_X1 port map( A => n11518, Z => n11392);
   U12366 : BUF_X1 port map( A => n11518, Z => n11391);
   U12367 : BUF_X1 port map( A => n11518, Z => n11390);
   U12368 : BUF_X1 port map( A => n11518, Z => n11389);
   U12369 : BUF_X1 port map( A => n11518, Z => n11394);
   U12370 : BUF_X1 port map( A => n11518, Z => n11399);
   U12371 : BUF_X1 port map( A => n11523, Z => n11340);
   U12372 : BUF_X1 port map( A => n11516, Z => n11421);
   U12373 : BUF_X1 port map( A => n11509, Z => n11508);
   U12374 : BUF_X1 port map( A => n11852, Z => n11766);
   U12375 : BUF_X1 port map( A => n11852, Z => n11767);
   U12376 : BUF_X1 port map( A => n11851, Z => n11768);
   U12377 : BUF_X1 port map( A => n11851, Z => n11769);
   U12378 : BUF_X1 port map( A => n11851, Z => n11770);
   U12379 : BUF_X1 port map( A => n11851, Z => n11771);
   U12380 : BUF_X1 port map( A => n11851, Z => n11772);
   U12381 : BUF_X1 port map( A => n11850, Z => n11773);
   U12382 : BUF_X1 port map( A => n11850, Z => n11774);
   U12383 : BUF_X1 port map( A => n11850, Z => n11775);
   U12384 : BUF_X1 port map( A => n11850, Z => n11776);
   U12385 : BUF_X1 port map( A => n11850, Z => n11777);
   U12386 : BUF_X1 port map( A => n11849, Z => n11778);
   U12387 : BUF_X1 port map( A => n11849, Z => n11779);
   U12388 : BUF_X1 port map( A => n11849, Z => n11780);
   U12389 : BUF_X1 port map( A => n11849, Z => n11781);
   U12390 : BUF_X1 port map( A => n11849, Z => n11782);
   U12391 : BUF_X1 port map( A => n11848, Z => n11783);
   U12392 : BUF_X1 port map( A => n11848, Z => n11784);
   U12393 : BUF_X1 port map( A => n11848, Z => n11785);
   U12394 : BUF_X1 port map( A => n11848, Z => n11786);
   U12395 : BUF_X1 port map( A => n11848, Z => n11787);
   U12396 : BUF_X1 port map( A => n11847, Z => n11788);
   U12397 : BUF_X1 port map( A => n11847, Z => n11789);
   U12398 : BUF_X1 port map( A => n11847, Z => n11790);
   U12399 : BUF_X1 port map( A => n11847, Z => n11791);
   U12400 : BUF_X1 port map( A => n11847, Z => n11792);
   U12401 : BUF_X1 port map( A => n11846, Z => n11793);
   U12402 : BUF_X1 port map( A => n11846, Z => n11794);
   U12403 : BUF_X1 port map( A => n11846, Z => n11795);
   U12404 : BUF_X1 port map( A => n11846, Z => n11796);
   U12405 : BUF_X1 port map( A => n11846, Z => n11797);
   U12406 : BUF_X1 port map( A => n11845, Z => n11798);
   U12407 : BUF_X1 port map( A => n11845, Z => n11799);
   U12408 : BUF_X1 port map( A => n11845, Z => n11800);
   U12409 : BUF_X1 port map( A => n11845, Z => n11801);
   U12410 : BUF_X1 port map( A => n11845, Z => n11802);
   U12411 : BUF_X1 port map( A => n11844, Z => n11803);
   U12412 : BUF_X1 port map( A => n11844, Z => n11804);
   U12413 : BUF_X1 port map( A => n11844, Z => n11805);
   U12414 : BUF_X1 port map( A => n11844, Z => n11806);
   U12415 : BUF_X1 port map( A => n11844, Z => n11807);
   U12416 : BUF_X1 port map( A => n11843, Z => n11808);
   U12417 : BUF_X1 port map( A => n11843, Z => n11809);
   U12418 : BUF_X1 port map( A => n11843, Z => n11810);
   U12419 : BUF_X1 port map( A => n11843, Z => n11811);
   U12420 : BUF_X1 port map( A => n11843, Z => n11812);
   U12421 : BUF_X1 port map( A => n11842, Z => n11813);
   U12422 : BUF_X1 port map( A => n11842, Z => n11814);
   U12423 : BUF_X1 port map( A => n11842, Z => n11815);
   U12424 : BUF_X1 port map( A => n11842, Z => n11816);
   U12425 : BUF_X1 port map( A => n11842, Z => n11817);
   U12426 : BUF_X1 port map( A => n11841, Z => n11818);
   U12427 : BUF_X1 port map( A => n11841, Z => n11819);
   U12428 : BUF_X1 port map( A => n11841, Z => n11820);
   U12429 : BUF_X1 port map( A => n11841, Z => n11821);
   U12430 : BUF_X1 port map( A => n11841, Z => n11822);
   U12431 : BUF_X1 port map( A => n11840, Z => n11823);
   U12432 : BUF_X1 port map( A => n11840, Z => n11824);
   U12433 : BUF_X1 port map( A => n11840, Z => n11825);
   U12434 : BUF_X1 port map( A => n11840, Z => n11826);
   U12435 : BUF_X1 port map( A => n11840, Z => n11827);
   U12436 : BUF_X1 port map( A => n11839, Z => n11828);
   U12437 : BUF_X1 port map( A => n11839, Z => n11829);
   U12438 : BUF_X1 port map( A => n11839, Z => n11830);
   U12439 : BUF_X1 port map( A => n11839, Z => n11831);
   U12440 : BUF_X1 port map( A => n11839, Z => n11832);
   U12441 : BUF_X1 port map( A => n11838, Z => n11833);
   U12442 : BUF_X1 port map( A => n11838, Z => n11834);
   U12443 : BUF_X1 port map( A => n11838, Z => n11835);
   U12444 : BUF_X1 port map( A => n11838, Z => n11836);
   U12445 : BUF_X1 port map( A => n11867, Z => n11688);
   U12446 : BUF_X1 port map( A => n11867, Z => n11689);
   U12447 : BUF_X1 port map( A => n11867, Z => n11690);
   U12448 : BUF_X1 port map( A => n11867, Z => n11691);
   U12449 : BUF_X1 port map( A => n11867, Z => n11692);
   U12450 : BUF_X1 port map( A => n11866, Z => n11693);
   U12451 : BUF_X1 port map( A => n11866, Z => n11694);
   U12452 : BUF_X1 port map( A => n11866, Z => n11695);
   U12453 : BUF_X1 port map( A => n11866, Z => n11696);
   U12454 : BUF_X1 port map( A => n11866, Z => n11697);
   U12455 : BUF_X1 port map( A => n11865, Z => n11698);
   U12456 : BUF_X1 port map( A => n11865, Z => n11699);
   U12457 : BUF_X1 port map( A => n11865, Z => n11700);
   U12458 : BUF_X1 port map( A => n11865, Z => n11701);
   U12459 : BUF_X1 port map( A => n11865, Z => n11702);
   U12460 : BUF_X1 port map( A => n11864, Z => n11703);
   U12461 : BUF_X1 port map( A => n11864, Z => n11704);
   U12462 : BUF_X1 port map( A => n11864, Z => n11705);
   U12463 : BUF_X1 port map( A => n11864, Z => n11706);
   U12464 : BUF_X1 port map( A => n11864, Z => n11707);
   U12465 : BUF_X1 port map( A => n11863, Z => n11708);
   U12466 : BUF_X1 port map( A => n11863, Z => n11709);
   U12467 : BUF_X1 port map( A => n11863, Z => n11710);
   U12468 : BUF_X1 port map( A => n11863, Z => n11711);
   U12469 : BUF_X1 port map( A => n11863, Z => n11712);
   U12470 : BUF_X1 port map( A => n11862, Z => n11713);
   U12471 : BUF_X1 port map( A => n11862, Z => n11714);
   U12472 : BUF_X1 port map( A => n11862, Z => n11715);
   U12473 : BUF_X1 port map( A => n11862, Z => n11716);
   U12474 : BUF_X1 port map( A => n11862, Z => n11717);
   U12475 : BUF_X1 port map( A => n11861, Z => n11718);
   U12476 : BUF_X1 port map( A => n11861, Z => n11719);
   U12477 : BUF_X1 port map( A => n11861, Z => n11720);
   U12478 : BUF_X1 port map( A => n11861, Z => n11721);
   U12479 : BUF_X1 port map( A => n11861, Z => n11722);
   U12480 : BUF_X1 port map( A => n11860, Z => n11723);
   U12481 : BUF_X1 port map( A => n11860, Z => n11724);
   U12482 : BUF_X1 port map( A => n11860, Z => n11725);
   U12483 : BUF_X1 port map( A => n11860, Z => n11726);
   U12484 : BUF_X1 port map( A => n11860, Z => n11727);
   U12485 : BUF_X1 port map( A => n11859, Z => n11728);
   U12486 : BUF_X1 port map( A => n11859, Z => n11729);
   U12487 : BUF_X1 port map( A => n11859, Z => n11730);
   U12488 : BUF_X1 port map( A => n11859, Z => n11731);
   U12489 : BUF_X1 port map( A => n11859, Z => n11732);
   U12490 : BUF_X1 port map( A => n11858, Z => n11733);
   U12491 : BUF_X1 port map( A => n11858, Z => n11734);
   U12492 : BUF_X1 port map( A => n11858, Z => n11735);
   U12493 : BUF_X1 port map( A => n11858, Z => n11736);
   U12494 : BUF_X1 port map( A => n11858, Z => n11737);
   U12495 : BUF_X1 port map( A => n11857, Z => n11738);
   U12496 : BUF_X1 port map( A => n11857, Z => n11739);
   U12497 : BUF_X1 port map( A => n11857, Z => n11740);
   U12498 : BUF_X1 port map( A => n11857, Z => n11741);
   U12499 : BUF_X1 port map( A => n11857, Z => n11742);
   U12500 : BUF_X1 port map( A => n11856, Z => n11743);
   U12501 : BUF_X1 port map( A => n11856, Z => n11744);
   U12502 : BUF_X1 port map( A => n11856, Z => n11745);
   U12503 : BUF_X1 port map( A => n11856, Z => n11746);
   U12504 : BUF_X1 port map( A => n11856, Z => n11747);
   U12505 : BUF_X1 port map( A => n11855, Z => n11748);
   U12506 : BUF_X1 port map( A => n11855, Z => n11749);
   U12507 : BUF_X1 port map( A => n11855, Z => n11750);
   U12508 : BUF_X1 port map( A => n11855, Z => n11751);
   U12509 : BUF_X1 port map( A => n11855, Z => n11752);
   U12510 : BUF_X1 port map( A => n11854, Z => n11753);
   U12511 : BUF_X1 port map( A => n11854, Z => n11754);
   U12512 : BUF_X1 port map( A => n11854, Z => n11755);
   U12513 : BUF_X1 port map( A => n11854, Z => n11756);
   U12514 : BUF_X1 port map( A => n11854, Z => n11757);
   U12515 : BUF_X1 port map( A => n11853, Z => n11758);
   U12516 : BUF_X1 port map( A => n11853, Z => n11759);
   U12517 : BUF_X1 port map( A => n11853, Z => n11760);
   U12518 : BUF_X1 port map( A => n11853, Z => n11761);
   U12519 : BUF_X1 port map( A => n11853, Z => n11762);
   U12520 : BUF_X1 port map( A => n11852, Z => n11763);
   U12521 : BUF_X1 port map( A => n11852, Z => n11764);
   U12522 : BUF_X1 port map( A => n11852, Z => n11765);
   U12523 : BUF_X1 port map( A => n11838, Z => n11837);
   U12524 : BUF_X1 port map( A => n11024, Z => n11013);
   U12525 : BUF_X1 port map( A => n11024, Z => n11014);
   U12526 : BUF_X1 port map( A => n11024, Z => n11015);
   U12527 : BUF_X1 port map( A => n11023, Z => n11016);
   U12528 : BUF_X1 port map( A => n11023, Z => n11017);
   U12529 : BUF_X1 port map( A => n11023, Z => n11018);
   U12530 : BUF_X1 port map( A => n10799, Z => n10788);
   U12531 : BUF_X1 port map( A => n10799, Z => n10789);
   U12532 : BUF_X1 port map( A => n10799, Z => n10790);
   U12533 : BUF_X1 port map( A => n10798, Z => n10791);
   U12534 : BUF_X1 port map( A => n10798, Z => n10792);
   U12535 : BUF_X1 port map( A => n10798, Z => n10793);
   U12536 : BUF_X1 port map( A => n11544, Z => n11542);
   U12537 : BUF_X1 port map( A => n11595, Z => n11593);
   U12538 : BUF_X1 port map( A => n11544, Z => n11541);
   U12539 : BUF_X1 port map( A => n11595, Z => n11592);
   U12540 : BUF_X1 port map( A => n11545, Z => n11540);
   U12541 : BUF_X1 port map( A => n11596, Z => n11591);
   U12542 : BUF_X1 port map( A => n11545, Z => n11539);
   U12543 : BUF_X1 port map( A => n11596, Z => n11590);
   U12544 : BUF_X1 port map( A => n11545, Z => n11538);
   U12545 : BUF_X1 port map( A => n11596, Z => n11589);
   U12546 : BUF_X1 port map( A => n11546, Z => n11537);
   U12547 : BUF_X1 port map( A => n11597, Z => n11588);
   U12548 : BUF_X1 port map( A => n11546, Z => n11536);
   U12549 : BUF_X1 port map( A => n11597, Z => n11587);
   U12550 : BUF_X1 port map( A => n11546, Z => n11535);
   U12551 : BUF_X1 port map( A => n11597, Z => n11586);
   U12552 : BUF_X1 port map( A => n11612, Z => n11610);
   U12553 : BUF_X1 port map( A => n11663, Z => n11661);
   U12554 : BUF_X1 port map( A => n11612, Z => n11609);
   U12555 : BUF_X1 port map( A => n11663, Z => n11660);
   U12556 : BUF_X1 port map( A => n11613, Z => n11608);
   U12557 : BUF_X1 port map( A => n11664, Z => n11659);
   U12558 : BUF_X1 port map( A => n11613, Z => n11607);
   U12559 : BUF_X1 port map( A => n11664, Z => n11658);
   U12560 : BUF_X1 port map( A => n11613, Z => n11606);
   U12561 : BUF_X1 port map( A => n11664, Z => n11657);
   U12562 : BUF_X1 port map( A => n11614, Z => n11605);
   U12563 : BUF_X1 port map( A => n11665, Z => n11656);
   U12564 : BUF_X1 port map( A => n11614, Z => n11604);
   U12565 : BUF_X1 port map( A => n11665, Z => n11655);
   U12566 : BUF_X1 port map( A => n11614, Z => n11603);
   U12567 : BUF_X1 port map( A => n11665, Z => n11654);
   U12568 : BUF_X1 port map( A => n10984, Z => n10982);
   U12569 : BUF_X1 port map( A => n10984, Z => n10981);
   U12570 : BUF_X1 port map( A => n10985, Z => n10980);
   U12571 : BUF_X1 port map( A => n10985, Z => n10979);
   U12572 : BUF_X1 port map( A => n10985, Z => n10978);
   U12573 : BUF_X1 port map( A => n10759, Z => n10757);
   U12574 : BUF_X1 port map( A => n10759, Z => n10756);
   U12575 : BUF_X1 port map( A => n10760, Z => n10755);
   U12576 : BUF_X1 port map( A => n10760, Z => n10754);
   U12577 : BUF_X1 port map( A => n10760, Z => n10753);
   U12578 : BUF_X1 port map( A => n11561, Z => n11559);
   U12579 : BUF_X1 port map( A => n11578, Z => n11576);
   U12580 : BUF_X1 port map( A => n11561, Z => n11558);
   U12581 : BUF_X1 port map( A => n11578, Z => n11575);
   U12582 : BUF_X1 port map( A => n11562, Z => n11557);
   U12583 : BUF_X1 port map( A => n11579, Z => n11574);
   U12584 : BUF_X1 port map( A => n11562, Z => n11556);
   U12585 : BUF_X1 port map( A => n11579, Z => n11573);
   U12586 : BUF_X1 port map( A => n11562, Z => n11555);
   U12587 : BUF_X1 port map( A => n11579, Z => n11572);
   U12588 : BUF_X1 port map( A => n11563, Z => n11554);
   U12589 : BUF_X1 port map( A => n11580, Z => n11571);
   U12590 : BUF_X1 port map( A => n11563, Z => n11553);
   U12591 : BUF_X1 port map( A => n11580, Z => n11570);
   U12592 : BUF_X1 port map( A => n11563, Z => n11552);
   U12593 : BUF_X1 port map( A => n11580, Z => n11569);
   U12594 : BUF_X1 port map( A => n11629, Z => n11627);
   U12595 : BUF_X1 port map( A => n11646, Z => n11644);
   U12596 : BUF_X1 port map( A => n11629, Z => n11626);
   U12597 : BUF_X1 port map( A => n11646, Z => n11643);
   U12598 : BUF_X1 port map( A => n11630, Z => n11625);
   U12599 : BUF_X1 port map( A => n11647, Z => n11642);
   U12600 : BUF_X1 port map( A => n11630, Z => n11624);
   U12601 : BUF_X1 port map( A => n11647, Z => n11641);
   U12602 : BUF_X1 port map( A => n11630, Z => n11623);
   U12603 : BUF_X1 port map( A => n11647, Z => n11640);
   U12604 : BUF_X1 port map( A => n11631, Z => n11622);
   U12605 : BUF_X1 port map( A => n11648, Z => n11639);
   U12606 : BUF_X1 port map( A => n11631, Z => n11621);
   U12607 : BUF_X1 port map( A => n11648, Z => n11638);
   U12608 : BUF_X1 port map( A => n11631, Z => n11620);
   U12609 : BUF_X1 port map( A => n11648, Z => n11637);
   U12610 : BUF_X1 port map( A => n10957, Z => n10955);
   U12611 : BUF_X1 port map( A => n10957, Z => n10954);
   U12612 : BUF_X1 port map( A => n10958, Z => n10953);
   U12613 : BUF_X1 port map( A => n10958, Z => n10952);
   U12614 : BUF_X1 port map( A => n10958, Z => n10951);
   U12615 : BUF_X1 port map( A => n10732, Z => n10730);
   U12616 : BUF_X1 port map( A => n10732, Z => n10729);
   U12617 : BUF_X1 port map( A => n10733, Z => n10728);
   U12618 : BUF_X1 port map( A => n10733, Z => n10727);
   U12619 : BUF_X1 port map( A => n10733, Z => n10726);
   U12620 : BUF_X1 port map( A => n10873, Z => n10871);
   U12621 : BUF_X1 port map( A => n10873, Z => n10870);
   U12622 : BUF_X1 port map( A => n10874, Z => n10869);
   U12623 : BUF_X1 port map( A => n10874, Z => n10868);
   U12624 : BUF_X1 port map( A => n10874, Z => n10867);
   U12625 : BUF_X1 port map( A => n10648, Z => n10646);
   U12626 : BUF_X1 port map( A => n10648, Z => n10645);
   U12627 : BUF_X1 port map( A => n10649, Z => n10644);
   U12628 : BUF_X1 port map( A => n10649, Z => n10643);
   U12629 : BUF_X1 port map( A => n10649, Z => n10642);
   U12630 : BUF_X1 port map( A => n10932, Z => n10930);
   U12631 : BUF_X1 port map( A => n10932, Z => n10929);
   U12632 : BUF_X1 port map( A => n10933, Z => n10928);
   U12633 : BUF_X1 port map( A => n10933, Z => n10927);
   U12634 : BUF_X1 port map( A => n10933, Z => n10926);
   U12635 : BUF_X1 port map( A => n10707, Z => n10705);
   U12636 : BUF_X1 port map( A => n10707, Z => n10704);
   U12637 : BUF_X1 port map( A => n10708, Z => n10703);
   U12638 : BUF_X1 port map( A => n10708, Z => n10702);
   U12639 : BUF_X1 port map( A => n10708, Z => n10701);
   U12640 : BUF_X1 port map( A => n11544, Z => n11543);
   U12641 : BUF_X1 port map( A => n11595, Z => n11594);
   U12642 : BUF_X1 port map( A => n11612, Z => n11611);
   U12643 : BUF_X1 port map( A => n11663, Z => n11662);
   U12644 : BUF_X1 port map( A => n11561, Z => n11560);
   U12645 : BUF_X1 port map( A => n11578, Z => n11577);
   U12646 : BUF_X1 port map( A => n11629, Z => n11628);
   U12647 : BUF_X1 port map( A => n11646, Z => n11645);
   U12648 : BUF_X1 port map( A => n11889, Z => n11887);
   U12649 : BUF_X1 port map( A => n11889, Z => n11886);
   U12650 : BUF_X1 port map( A => n11890, Z => n11885);
   U12651 : BUF_X1 port map( A => n11890, Z => n11884);
   U12652 : BUF_X1 port map( A => n11890, Z => n11883);
   U12653 : BUF_X1 port map( A => n10984, Z => n10983);
   U12654 : BUF_X1 port map( A => n10759, Z => n10758);
   U12655 : BUF_X1 port map( A => n10957, Z => n10956);
   U12656 : BUF_X1 port map( A => n10732, Z => n10731);
   U12657 : BUF_X1 port map( A => n10873, Z => n10872);
   U12658 : BUF_X1 port map( A => n10648, Z => n10647);
   U12659 : BUF_X1 port map( A => n10932, Z => n10931);
   U12660 : BUF_X1 port map( A => n10707, Z => n10706);
   U12661 : BUF_X1 port map( A => n11889, Z => n11888);
   U12662 : BUF_X1 port map( A => n11871, Z => n11668);
   U12663 : BUF_X1 port map( A => n11871, Z => n11669);
   U12664 : BUF_X1 port map( A => n11871, Z => n11670);
   U12665 : BUF_X1 port map( A => n11871, Z => n11671);
   U12666 : BUF_X1 port map( A => n11871, Z => n11672);
   U12667 : BUF_X1 port map( A => n11870, Z => n11673);
   U12668 : BUF_X1 port map( A => n11870, Z => n11674);
   U12669 : BUF_X1 port map( A => n11870, Z => n11675);
   U12670 : BUF_X1 port map( A => n11870, Z => n11676);
   U12671 : BUF_X1 port map( A => n11870, Z => n11677);
   U12672 : BUF_X1 port map( A => n11869, Z => n11678);
   U12673 : BUF_X1 port map( A => n11869, Z => n11679);
   U12674 : BUF_X1 port map( A => n11869, Z => n11680);
   U12675 : BUF_X1 port map( A => n11869, Z => n11681);
   U12676 : BUF_X1 port map( A => n11869, Z => n11682);
   U12677 : BUF_X1 port map( A => n11868, Z => n11683);
   U12678 : BUF_X1 port map( A => n11868, Z => n11684);
   U12679 : BUF_X1 port map( A => n11868, Z => n11685);
   U12680 : BUF_X1 port map( A => n11868, Z => n11686);
   U12681 : BUF_X1 port map( A => n11868, Z => n11687);
   U12682 : BUF_X1 port map( A => n11877, Z => n11851);
   U12683 : BUF_X1 port map( A => n11877, Z => n11850);
   U12684 : BUF_X1 port map( A => n11877, Z => n11849);
   U12685 : BUF_X1 port map( A => n11877, Z => n11848);
   U12686 : BUF_X1 port map( A => n11878, Z => n11847);
   U12687 : BUF_X1 port map( A => n11878, Z => n11846);
   U12688 : BUF_X1 port map( A => n11878, Z => n11845);
   U12689 : BUF_X1 port map( A => n11878, Z => n11844);
   U12690 : BUF_X1 port map( A => n11878, Z => n11843);
   U12691 : BUF_X1 port map( A => n11879, Z => n11842);
   U12692 : BUF_X1 port map( A => n11879, Z => n11841);
   U12693 : BUF_X1 port map( A => n11879, Z => n11840);
   U12694 : BUF_X1 port map( A => n11879, Z => n11839);
   U12695 : BUF_X1 port map( A => n11879, Z => n11838);
   U12696 : BUF_X1 port map( A => n11874, Z => n11867);
   U12697 : BUF_X1 port map( A => n11874, Z => n11866);
   U12698 : BUF_X1 port map( A => n11874, Z => n11865);
   U12699 : BUF_X1 port map( A => n11874, Z => n11864);
   U12700 : BUF_X1 port map( A => n11874, Z => n11863);
   U12701 : BUF_X1 port map( A => n11875, Z => n11862);
   U12702 : BUF_X1 port map( A => n11875, Z => n11861);
   U12703 : BUF_X1 port map( A => n11875, Z => n11860);
   U12704 : BUF_X1 port map( A => n11875, Z => n11859);
   U12705 : BUF_X1 port map( A => n11875, Z => n11858);
   U12706 : BUF_X1 port map( A => n11876, Z => n11857);
   U12707 : BUF_X1 port map( A => n11876, Z => n11856);
   U12708 : BUF_X1 port map( A => n11876, Z => n11855);
   U12709 : BUF_X1 port map( A => n11876, Z => n11854);
   U12710 : BUF_X1 port map( A => n11876, Z => n11853);
   U12711 : BUF_X1 port map( A => n11877, Z => n11852);
   U12712 : BUF_X1 port map( A => n11022, Z => n11019);
   U12713 : BUF_X1 port map( A => n11022, Z => n11020);
   U12714 : BUF_X1 port map( A => n10797, Z => n10794);
   U12715 : BUF_X1 port map( A => n10797, Z => n10795);
   U12716 : BUF_X1 port map( A => n11025, Z => n11012);
   U12717 : BUF_X1 port map( A => n11026, Z => n11025);
   U12718 : BUF_X1 port map( A => n10800, Z => n10787);
   U12719 : BUF_X1 port map( A => n10801, Z => n10800);
   U12720 : BUF_X1 port map( A => n11007, Z => n10996);
   U12721 : BUF_X1 port map( A => n11007, Z => n10997);
   U12722 : BUF_X1 port map( A => n11007, Z => n10998);
   U12723 : BUF_X1 port map( A => n11006, Z => n10999);
   U12724 : BUF_X1 port map( A => n11006, Z => n11000);
   U12725 : BUF_X1 port map( A => n11006, Z => n11001);
   U12726 : BUF_X1 port map( A => n10782, Z => n10771);
   U12727 : BUF_X1 port map( A => n10782, Z => n10772);
   U12728 : BUF_X1 port map( A => n10782, Z => n10773);
   U12729 : BUF_X1 port map( A => n10781, Z => n10774);
   U12730 : BUF_X1 port map( A => n10781, Z => n10775);
   U12731 : BUF_X1 port map( A => n10781, Z => n10776);
   U12732 : BUF_X1 port map( A => n11022, Z => n11021);
   U12733 : BUF_X1 port map( A => n10797, Z => n10796);
   U12734 : BUF_X1 port map( A => n10865, Z => n10863);
   U12735 : BUF_X1 port map( A => n10865, Z => n10862);
   U12736 : BUF_X1 port map( A => n10866, Z => n10861);
   U12737 : BUF_X1 port map( A => n10866, Z => n10860);
   U12738 : BUF_X1 port map( A => n10866, Z => n10859);
   U12739 : BUF_X1 port map( A => n10640, Z => n10638);
   U12740 : BUF_X1 port map( A => n10640, Z => n10637);
   U12741 : BUF_X1 port map( A => n10641, Z => n10636);
   U12742 : BUF_X1 port map( A => n10641, Z => n10635);
   U12743 : BUF_X1 port map( A => n10641, Z => n10634);
   U12744 : BUF_X1 port map( A => n11547, Z => n11534);
   U12745 : BUF_X1 port map( A => n11598, Z => n11585);
   U12746 : BUF_X1 port map( A => n11547, Z => n11533);
   U12747 : BUF_X1 port map( A => n11598, Z => n11584);
   U12748 : BUF_X1 port map( A => n11615, Z => n11602);
   U12749 : BUF_X1 port map( A => n11666, Z => n11653);
   U12750 : BUF_X1 port map( A => n11615, Z => n11601);
   U12751 : BUF_X1 port map( A => n11666, Z => n11652);
   U12752 : BUF_X1 port map( A => n10856, Z => n10854);
   U12753 : BUF_X1 port map( A => n10975, Z => n10973);
   U12754 : BUF_X1 port map( A => n10856, Z => n10853);
   U12755 : BUF_X1 port map( A => n10975, Z => n10972);
   U12756 : BUF_X1 port map( A => n10857, Z => n10852);
   U12757 : BUF_X1 port map( A => n10976, Z => n10971);
   U12758 : BUF_X1 port map( A => n10857, Z => n10851);
   U12759 : BUF_X1 port map( A => n10976, Z => n10970);
   U12760 : BUF_X1 port map( A => n10857, Z => n10850);
   U12761 : BUF_X1 port map( A => n10976, Z => n10969);
   U12762 : BUF_X1 port map( A => n10631, Z => n10629);
   U12763 : BUF_X1 port map( A => n10750, Z => n10748);
   U12764 : BUF_X1 port map( A => n10631, Z => n10628);
   U12765 : BUF_X1 port map( A => n10750, Z => n10747);
   U12766 : BUF_X1 port map( A => n10632, Z => n10627);
   U12767 : BUF_X1 port map( A => n10751, Z => n10746);
   U12768 : BUF_X1 port map( A => n10632, Z => n10626);
   U12769 : BUF_X1 port map( A => n10751, Z => n10745);
   U12770 : BUF_X1 port map( A => n10632, Z => n10625);
   U12771 : BUF_X1 port map( A => n10751, Z => n10744);
   U12772 : BUF_X1 port map( A => n11564, Z => n11551);
   U12773 : BUF_X1 port map( A => n11581, Z => n11568);
   U12774 : BUF_X1 port map( A => n11564, Z => n11550);
   U12775 : BUF_X1 port map( A => n11581, Z => n11567);
   U12776 : BUF_X1 port map( A => n11632, Z => n11619);
   U12777 : BUF_X1 port map( A => n11649, Z => n11636);
   U12778 : BUF_X1 port map( A => n11632, Z => n11618);
   U12779 : BUF_X1 port map( A => n11649, Z => n11635);
   U12780 : BUF_X1 port map( A => n11060, Z => n11049);
   U12781 : BUF_X1 port map( A => n11060, Z => n11050);
   U12782 : BUF_X1 port map( A => n11060, Z => n11051);
   U12783 : BUF_X1 port map( A => n11059, Z => n11052);
   U12784 : BUF_X1 port map( A => n11059, Z => n11053);
   U12785 : BUF_X1 port map( A => n11059, Z => n11054);
   U12786 : BUF_X1 port map( A => n10835, Z => n10824);
   U12787 : BUF_X1 port map( A => n10835, Z => n10825);
   U12788 : BUF_X1 port map( A => n10835, Z => n10826);
   U12789 : BUF_X1 port map( A => n10834, Z => n10827);
   U12790 : BUF_X1 port map( A => n10834, Z => n10828);
   U12791 : BUF_X1 port map( A => n10834, Z => n10829);
   U12792 : BUF_X1 port map( A => n10924, Z => n10922);
   U12793 : BUF_X1 port map( A => n10881, Z => n10879);
   U12794 : BUF_X1 port map( A => n10924, Z => n10921);
   U12795 : BUF_X1 port map( A => n10881, Z => n10878);
   U12796 : BUF_X1 port map( A => n10925, Z => n10920);
   U12797 : BUF_X1 port map( A => n10882, Z => n10877);
   U12798 : BUF_X1 port map( A => n10925, Z => n10919);
   U12799 : BUF_X1 port map( A => n10882, Z => n10876);
   U12800 : BUF_X1 port map( A => n10925, Z => n10918);
   U12801 : BUF_X1 port map( A => n10882, Z => n10875);
   U12802 : BUF_X1 port map( A => n10699, Z => n10697);
   U12803 : BUF_X1 port map( A => n10656, Z => n10654);
   U12804 : BUF_X1 port map( A => n10699, Z => n10696);
   U12805 : BUF_X1 port map( A => n10656, Z => n10653);
   U12806 : BUF_X1 port map( A => n10700, Z => n10695);
   U12807 : BUF_X1 port map( A => n10657, Z => n10652);
   U12808 : BUF_X1 port map( A => n10700, Z => n10694);
   U12809 : BUF_X1 port map( A => n10657, Z => n10651);
   U12810 : BUF_X1 port map( A => n10700, Z => n10693);
   U12811 : BUF_X1 port map( A => n10657, Z => n10650);
   U12812 : BUF_X1 port map( A => n11061, Z => n11047);
   U12813 : BUF_X1 port map( A => n11061, Z => n11048);
   U12814 : BUF_X1 port map( A => n10836, Z => n10822);
   U12815 : BUF_X1 port map( A => n10836, Z => n10823);
   U12816 : BUF_X1 port map( A => n10948, Z => n10946);
   U12817 : BUF_X1 port map( A => n10948, Z => n10945);
   U12818 : BUF_X1 port map( A => n10949, Z => n10944);
   U12819 : BUF_X1 port map( A => n10949, Z => n10943);
   U12820 : BUF_X1 port map( A => n10949, Z => n10942);
   U12821 : BUF_X1 port map( A => n10723, Z => n10721);
   U12822 : BUF_X1 port map( A => n10723, Z => n10720);
   U12823 : BUF_X1 port map( A => n10724, Z => n10719);
   U12824 : BUF_X1 port map( A => n10724, Z => n10718);
   U12825 : BUF_X1 port map( A => n10724, Z => n10717);
   U12826 : BUF_X1 port map( A => n11042, Z => n11031);
   U12827 : BUF_X1 port map( A => n11042, Z => n11032);
   U12828 : BUF_X1 port map( A => n11042, Z => n11033);
   U12829 : BUF_X1 port map( A => n11041, Z => n11034);
   U12830 : BUF_X1 port map( A => n11041, Z => n11035);
   U12831 : BUF_X1 port map( A => n11041, Z => n11036);
   U12832 : BUF_X1 port map( A => n10817, Z => n10806);
   U12833 : BUF_X1 port map( A => n10817, Z => n10807);
   U12834 : BUF_X1 port map( A => n10817, Z => n10808);
   U12835 : BUF_X1 port map( A => n10816, Z => n10809);
   U12836 : BUF_X1 port map( A => n10816, Z => n10810);
   U12837 : BUF_X1 port map( A => n10816, Z => n10811);
   U12838 : BUF_X1 port map( A => n10916, Z => n10914);
   U12839 : BUF_X1 port map( A => n10916, Z => n10913);
   U12840 : BUF_X1 port map( A => n10917, Z => n10912);
   U12841 : BUF_X1 port map( A => n10917, Z => n10911);
   U12842 : BUF_X1 port map( A => n10917, Z => n10910);
   U12843 : BUF_X1 port map( A => n10691, Z => n10689);
   U12844 : BUF_X1 port map( A => n10691, Z => n10688);
   U12845 : BUF_X1 port map( A => n10692, Z => n10687);
   U12846 : BUF_X1 port map( A => n10692, Z => n10686);
   U12847 : BUF_X1 port map( A => n10692, Z => n10685);
   U12848 : BUF_X1 port map( A => n11072, Z => n11070);
   U12849 : BUF_X1 port map( A => n11072, Z => n11069);
   U12850 : BUF_X1 port map( A => n11073, Z => n11068);
   U12851 : BUF_X1 port map( A => n11073, Z => n11067);
   U12852 : BUF_X1 port map( A => n11073, Z => n11066);
   U12853 : BUF_X1 port map( A => n10847, Z => n10845);
   U12854 : BUF_X1 port map( A => n10847, Z => n10844);
   U12855 : BUF_X1 port map( A => n10848, Z => n10843);
   U12856 : BUF_X1 port map( A => n10848, Z => n10842);
   U12857 : BUF_X1 port map( A => n10848, Z => n10841);
   U12858 : BUF_X1 port map( A => n10966, Z => n10964);
   U12859 : BUF_X1 port map( A => n10966, Z => n10963);
   U12860 : BUF_X1 port map( A => n10967, Z => n10962);
   U12861 : BUF_X1 port map( A => n10967, Z => n10961);
   U12862 : BUF_X1 port map( A => n10967, Z => n10960);
   U12863 : BUF_X1 port map( A => n10741, Z => n10739);
   U12864 : BUF_X1 port map( A => n10741, Z => n10738);
   U12865 : BUF_X1 port map( A => n10742, Z => n10737);
   U12866 : BUF_X1 port map( A => n10742, Z => n10736);
   U12867 : BUF_X1 port map( A => n10742, Z => n10735);
   U12868 : BUF_X1 port map( A => n11043, Z => n11029);
   U12869 : BUF_X1 port map( A => n11043, Z => n11030);
   U12870 : BUF_X1 port map( A => n10818, Z => n10804);
   U12871 : BUF_X1 port map( A => n10818, Z => n10805);
   U12872 : BUF_X1 port map( A => n10890, Z => n10888);
   U12873 : BUF_X1 port map( A => n10890, Z => n10887);
   U12874 : BUF_X1 port map( A => n10891, Z => n10886);
   U12875 : BUF_X1 port map( A => n10891, Z => n10885);
   U12876 : BUF_X1 port map( A => n10891, Z => n10884);
   U12877 : BUF_X1 port map( A => n10665, Z => n10663);
   U12878 : BUF_X1 port map( A => n10665, Z => n10662);
   U12879 : BUF_X1 port map( A => n10666, Z => n10661);
   U12880 : BUF_X1 port map( A => n10666, Z => n10660);
   U12881 : BUF_X1 port map( A => n10666, Z => n10659);
   U12882 : BUF_X1 port map( A => n10940, Z => n10938);
   U12883 : BUF_X1 port map( A => n10940, Z => n10937);
   U12884 : BUF_X1 port map( A => n10941, Z => n10936);
   U12885 : BUF_X1 port map( A => n10941, Z => n10935);
   U12886 : BUF_X1 port map( A => n10941, Z => n10934);
   U12887 : BUF_X1 port map( A => n10715, Z => n10713);
   U12888 : BUF_X1 port map( A => n10715, Z => n10712);
   U12889 : BUF_X1 port map( A => n10716, Z => n10711);
   U12890 : BUF_X1 port map( A => n10716, Z => n10710);
   U12891 : BUF_X1 port map( A => n10716, Z => n10709);
   U12892 : BUF_X1 port map( A => n10899, Z => n10897);
   U12893 : BUF_X1 port map( A => n10899, Z => n10896);
   U12894 : BUF_X1 port map( A => n10900, Z => n10895);
   U12895 : BUF_X1 port map( A => n10900, Z => n10894);
   U12896 : BUF_X1 port map( A => n10900, Z => n10893);
   U12897 : BUF_X1 port map( A => n10674, Z => n10672);
   U12898 : BUF_X1 port map( A => n10674, Z => n10671);
   U12899 : BUF_X1 port map( A => n10675, Z => n10670);
   U12900 : BUF_X1 port map( A => n10675, Z => n10669);
   U12901 : BUF_X1 port map( A => n10675, Z => n10668);
   U12902 : BUF_X1 port map( A => n10908, Z => n10906);
   U12903 : BUF_X1 port map( A => n10908, Z => n10905);
   U12904 : BUF_X1 port map( A => n10909, Z => n10904);
   U12905 : BUF_X1 port map( A => n10909, Z => n10903);
   U12906 : BUF_X1 port map( A => n10909, Z => n10902);
   U12907 : BUF_X1 port map( A => n10683, Z => n10681);
   U12908 : BUF_X1 port map( A => n10683, Z => n10680);
   U12909 : BUF_X1 port map( A => n10684, Z => n10679);
   U12910 : BUF_X1 port map( A => n10684, Z => n10678);
   U12911 : BUF_X1 port map( A => n10684, Z => n10677);
   U12912 : BUF_X1 port map( A => n11527, Z => n11513);
   U12913 : BUF_X1 port map( A => n11526, Z => n11515);
   U12914 : BUF_X1 port map( A => n11527, Z => n11514);
   U12915 : BUF_X1 port map( A => n11528, Z => n11509);
   U12916 : BUF_X1 port map( A => n11527, Z => n11512);
   U12917 : BUF_X1 port map( A => n11528, Z => n11511);
   U12918 : BUF_X1 port map( A => n11528, Z => n11510);
   U12919 : BUF_X1 port map( A => n11525, Z => n11520);
   U12920 : BUF_X1 port map( A => n11524, Z => n11522);
   U12921 : BUF_X1 port map( A => n11524, Z => n11521);
   U12922 : BUF_X1 port map( A => n11526, Z => n11517);
   U12923 : BUF_X1 port map( A => n11525, Z => n11519);
   U12924 : BUF_X1 port map( A => n11525, Z => n11518);
   U12925 : BUF_X1 port map( A => n11526, Z => n11516);
   U12926 : BUF_X1 port map( A => n11524, Z => n11523);
   U12927 : BUF_X1 port map( A => n12169, Z => n12162);
   U12928 : BUF_X1 port map( A => n12169, Z => n12163);
   U12929 : BUF_X1 port map( A => n12169, Z => n12164);
   U12930 : BUF_X1 port map( A => n12168, Z => n12165);
   U12931 : BUF_X1 port map( A => n12168, Z => n12166);
   U12932 : BUF_X1 port map( A => n12160, Z => n12153);
   U12933 : BUF_X1 port map( A => n12160, Z => n12154);
   U12934 : BUF_X1 port map( A => n12160, Z => n12155);
   U12935 : BUF_X1 port map( A => n12159, Z => n12156);
   U12936 : BUF_X1 port map( A => n12159, Z => n12157);
   U12937 : BUF_X1 port map( A => n12150, Z => n12148);
   U12938 : BUF_X1 port map( A => n12150, Z => n12147);
   U12939 : BUF_X1 port map( A => n12151, Z => n12146);
   U12940 : BUF_X1 port map( A => n12151, Z => n12145);
   U12941 : BUF_X1 port map( A => n12151, Z => n12144);
   U12942 : BUF_X1 port map( A => n12141, Z => n12139);
   U12943 : BUF_X1 port map( A => n12141, Z => n12138);
   U12944 : BUF_X1 port map( A => n12142, Z => n12137);
   U12945 : BUF_X1 port map( A => n12142, Z => n12136);
   U12946 : BUF_X1 port map( A => n12142, Z => n12135);
   U12947 : BUF_X1 port map( A => n12132, Z => n12130);
   U12948 : BUF_X1 port map( A => n12132, Z => n12129);
   U12949 : BUF_X1 port map( A => n12133, Z => n12128);
   U12950 : BUF_X1 port map( A => n12133, Z => n12127);
   U12951 : BUF_X1 port map( A => n12133, Z => n12126);
   U12952 : BUF_X1 port map( A => n12123, Z => n12121);
   U12953 : BUF_X1 port map( A => n12123, Z => n12120);
   U12954 : BUF_X1 port map( A => n12124, Z => n12119);
   U12955 : BUF_X1 port map( A => n12124, Z => n12118);
   U12956 : BUF_X1 port map( A => n12124, Z => n12117);
   U12957 : BUF_X1 port map( A => n12114, Z => n12112);
   U12958 : BUF_X1 port map( A => n12114, Z => n12111);
   U12959 : BUF_X1 port map( A => n12115, Z => n12110);
   U12960 : BUF_X1 port map( A => n12115, Z => n12109);
   U12961 : BUF_X1 port map( A => n12115, Z => n12108);
   U12962 : BUF_X1 port map( A => n12105, Z => n12103);
   U12963 : BUF_X1 port map( A => n12105, Z => n12102);
   U12964 : BUF_X1 port map( A => n12106, Z => n12101);
   U12965 : BUF_X1 port map( A => n12106, Z => n12100);
   U12966 : BUF_X1 port map( A => n12106, Z => n12099);
   U12967 : BUF_X1 port map( A => n12096, Z => n12094);
   U12968 : BUF_X1 port map( A => n12096, Z => n12093);
   U12969 : BUF_X1 port map( A => n12097, Z => n12092);
   U12970 : BUF_X1 port map( A => n12097, Z => n12091);
   U12971 : BUF_X1 port map( A => n12097, Z => n12090);
   U12972 : BUF_X1 port map( A => n12087, Z => n12085);
   U12973 : BUF_X1 port map( A => n12087, Z => n12084);
   U12974 : BUF_X1 port map( A => n12088, Z => n12083);
   U12975 : BUF_X1 port map( A => n12088, Z => n12082);
   U12976 : BUF_X1 port map( A => n12088, Z => n12081);
   U12977 : BUF_X1 port map( A => n12078, Z => n12076);
   U12978 : BUF_X1 port map( A => n12078, Z => n12075);
   U12979 : BUF_X1 port map( A => n12079, Z => n12074);
   U12980 : BUF_X1 port map( A => n12079, Z => n12073);
   U12981 : BUF_X1 port map( A => n12079, Z => n12072);
   U12982 : BUF_X1 port map( A => n12069, Z => n12067);
   U12983 : BUF_X1 port map( A => n12069, Z => n12066);
   U12984 : BUF_X1 port map( A => n12070, Z => n12065);
   U12985 : BUF_X1 port map( A => n12070, Z => n12064);
   U12986 : BUF_X1 port map( A => n12070, Z => n12063);
   U12987 : BUF_X1 port map( A => n12060, Z => n12058);
   U12988 : BUF_X1 port map( A => n12060, Z => n12057);
   U12989 : BUF_X1 port map( A => n12061, Z => n12056);
   U12990 : BUF_X1 port map( A => n12061, Z => n12055);
   U12991 : BUF_X1 port map( A => n12061, Z => n12054);
   U12992 : BUF_X1 port map( A => n12051, Z => n12049);
   U12993 : BUF_X1 port map( A => n12051, Z => n12048);
   U12994 : BUF_X1 port map( A => n12052, Z => n12047);
   U12995 : BUF_X1 port map( A => n12052, Z => n12046);
   U12996 : BUF_X1 port map( A => n12052, Z => n12045);
   U12997 : BUF_X1 port map( A => n12042, Z => n12040);
   U12998 : BUF_X1 port map( A => n12042, Z => n12039);
   U12999 : BUF_X1 port map( A => n12043, Z => n12038);
   U13000 : BUF_X1 port map( A => n12043, Z => n12037);
   U13001 : BUF_X1 port map( A => n12043, Z => n12036);
   U13002 : BUF_X1 port map( A => n12033, Z => n12031);
   U13003 : BUF_X1 port map( A => n12033, Z => n12030);
   U13004 : BUF_X1 port map( A => n12034, Z => n12029);
   U13005 : BUF_X1 port map( A => n12034, Z => n12028);
   U13006 : BUF_X1 port map( A => n12034, Z => n12027);
   U13007 : BUF_X1 port map( A => n12024, Z => n12022);
   U13008 : BUF_X1 port map( A => n12024, Z => n12021);
   U13009 : BUF_X1 port map( A => n12025, Z => n12020);
   U13010 : BUF_X1 port map( A => n12025, Z => n12019);
   U13011 : BUF_X1 port map( A => n12025, Z => n12018);
   U13012 : BUF_X1 port map( A => n12015, Z => n12013);
   U13013 : BUF_X1 port map( A => n12015, Z => n12012);
   U13014 : BUF_X1 port map( A => n12016, Z => n12011);
   U13015 : BUF_X1 port map( A => n12016, Z => n12010);
   U13016 : BUF_X1 port map( A => n12016, Z => n12009);
   U13017 : BUF_X1 port map( A => n12006, Z => n12004);
   U13018 : BUF_X1 port map( A => n12006, Z => n12003);
   U13019 : BUF_X1 port map( A => n12007, Z => n12002);
   U13020 : BUF_X1 port map( A => n12007, Z => n12001);
   U13021 : BUF_X1 port map( A => n12007, Z => n12000);
   U13022 : BUF_X1 port map( A => n11997, Z => n11995);
   U13023 : BUF_X1 port map( A => n11997, Z => n11994);
   U13024 : BUF_X1 port map( A => n11998, Z => n11993);
   U13025 : BUF_X1 port map( A => n11998, Z => n11992);
   U13026 : BUF_X1 port map( A => n11998, Z => n11991);
   U13027 : BUF_X1 port map( A => n11988, Z => n11986);
   U13028 : BUF_X1 port map( A => n11988, Z => n11985);
   U13029 : BUF_X1 port map( A => n11989, Z => n11984);
   U13030 : BUF_X1 port map( A => n11989, Z => n11983);
   U13031 : BUF_X1 port map( A => n11989, Z => n11982);
   U13032 : BUF_X1 port map( A => n11979, Z => n11977);
   U13033 : BUF_X1 port map( A => n11979, Z => n11976);
   U13034 : BUF_X1 port map( A => n11980, Z => n11975);
   U13035 : BUF_X1 port map( A => n11980, Z => n11974);
   U13036 : BUF_X1 port map( A => n11980, Z => n11973);
   U13037 : BUF_X1 port map( A => n11970, Z => n11968);
   U13038 : BUF_X1 port map( A => n11970, Z => n11967);
   U13039 : BUF_X1 port map( A => n11971, Z => n11966);
   U13040 : BUF_X1 port map( A => n11971, Z => n11965);
   U13041 : BUF_X1 port map( A => n11971, Z => n11964);
   U13042 : BUF_X1 port map( A => n11961, Z => n11959);
   U13043 : BUF_X1 port map( A => n11961, Z => n11958);
   U13044 : BUF_X1 port map( A => n11962, Z => n11957);
   U13045 : BUF_X1 port map( A => n11962, Z => n11956);
   U13046 : BUF_X1 port map( A => n11962, Z => n11955);
   U13047 : BUF_X1 port map( A => n11952, Z => n11950);
   U13048 : BUF_X1 port map( A => n11952, Z => n11949);
   U13049 : BUF_X1 port map( A => n11953, Z => n11948);
   U13050 : BUF_X1 port map( A => n11953, Z => n11947);
   U13051 : BUF_X1 port map( A => n11953, Z => n11946);
   U13052 : BUF_X1 port map( A => n11943, Z => n11941);
   U13053 : BUF_X1 port map( A => n11943, Z => n11940);
   U13054 : BUF_X1 port map( A => n11944, Z => n11939);
   U13055 : BUF_X1 port map( A => n11944, Z => n11938);
   U13056 : BUF_X1 port map( A => n11944, Z => n11937);
   U13057 : BUF_X1 port map( A => n11934, Z => n11932);
   U13058 : BUF_X1 port map( A => n11934, Z => n11931);
   U13059 : BUF_X1 port map( A => n11935, Z => n11930);
   U13060 : BUF_X1 port map( A => n11935, Z => n11929);
   U13061 : BUF_X1 port map( A => n11935, Z => n11928);
   U13062 : BUF_X1 port map( A => n11925, Z => n11923);
   U13063 : BUF_X1 port map( A => n11925, Z => n11922);
   U13064 : BUF_X1 port map( A => n11926, Z => n11921);
   U13065 : BUF_X1 port map( A => n11926, Z => n11920);
   U13066 : BUF_X1 port map( A => n11926, Z => n11919);
   U13067 : BUF_X1 port map( A => n11916, Z => n11914);
   U13068 : BUF_X1 port map( A => n11916, Z => n11913);
   U13069 : BUF_X1 port map( A => n11917, Z => n11912);
   U13070 : BUF_X1 port map( A => n11917, Z => n11911);
   U13071 : BUF_X1 port map( A => n11917, Z => n11910);
   U13072 : BUF_X1 port map( A => n11907, Z => n11905);
   U13073 : BUF_X1 port map( A => n11907, Z => n11904);
   U13074 : BUF_X1 port map( A => n11908, Z => n11903);
   U13075 : BUF_X1 port map( A => n11908, Z => n11902);
   U13076 : BUF_X1 port map( A => n11908, Z => n11901);
   U13077 : BUF_X1 port map( A => n11898, Z => n11896);
   U13078 : BUF_X1 port map( A => n11898, Z => n11895);
   U13079 : BUF_X1 port map( A => n11899, Z => n11894);
   U13080 : BUF_X1 port map( A => n11899, Z => n11893);
   U13081 : BUF_X1 port map( A => n11899, Z => n11892);
   U13082 : BUF_X1 port map( A => n10865, Z => n10864);
   U13083 : BUF_X1 port map( A => n10640, Z => n10639);
   U13084 : BUF_X1 port map( A => n10856, Z => n10855);
   U13085 : BUF_X1 port map( A => n10975, Z => n10974);
   U13086 : BUF_X1 port map( A => n10631, Z => n10630);
   U13087 : BUF_X1 port map( A => n10750, Z => n10749);
   U13088 : BUF_X1 port map( A => n10924, Z => n10923);
   U13089 : BUF_X1 port map( A => n10881, Z => n10880);
   U13090 : BUF_X1 port map( A => n10699, Z => n10698);
   U13091 : BUF_X1 port map( A => n10656, Z => n10655);
   U13092 : BUF_X1 port map( A => n10948, Z => n10947);
   U13093 : BUF_X1 port map( A => n10723, Z => n10722);
   U13094 : BUF_X1 port map( A => n10916, Z => n10915);
   U13095 : BUF_X1 port map( A => n10691, Z => n10690);
   U13096 : BUF_X1 port map( A => n11072, Z => n11071);
   U13097 : BUF_X1 port map( A => n10847, Z => n10846);
   U13098 : BUF_X1 port map( A => n10966, Z => n10965);
   U13099 : BUF_X1 port map( A => n10741, Z => n10740);
   U13100 : BUF_X1 port map( A => n10890, Z => n10889);
   U13101 : BUF_X1 port map( A => n10665, Z => n10664);
   U13102 : BUF_X1 port map( A => n10940, Z => n10939);
   U13103 : BUF_X1 port map( A => n10715, Z => n10714);
   U13104 : BUF_X1 port map( A => n10899, Z => n10898);
   U13105 : BUF_X1 port map( A => n10674, Z => n10673);
   U13106 : BUF_X1 port map( A => n10908, Z => n10907);
   U13107 : BUF_X1 port map( A => n10683, Z => n10682);
   U13108 : BUF_X1 port map( A => n12168, Z => n12167);
   U13109 : BUF_X1 port map( A => n12159, Z => n12158);
   U13110 : BUF_X1 port map( A => n12150, Z => n12149);
   U13111 : BUF_X1 port map( A => n12141, Z => n12140);
   U13112 : BUF_X1 port map( A => n12132, Z => n12131);
   U13113 : BUF_X1 port map( A => n12123, Z => n12122);
   U13114 : BUF_X1 port map( A => n12114, Z => n12113);
   U13115 : BUF_X1 port map( A => n12105, Z => n12104);
   U13116 : BUF_X1 port map( A => n12096, Z => n12095);
   U13117 : BUF_X1 port map( A => n12087, Z => n12086);
   U13118 : BUF_X1 port map( A => n12078, Z => n12077);
   U13119 : BUF_X1 port map( A => n12069, Z => n12068);
   U13120 : BUF_X1 port map( A => n12060, Z => n12059);
   U13121 : BUF_X1 port map( A => n12051, Z => n12050);
   U13122 : BUF_X1 port map( A => n12042, Z => n12041);
   U13123 : BUF_X1 port map( A => n12033, Z => n12032);
   U13124 : BUF_X1 port map( A => n12024, Z => n12023);
   U13125 : BUF_X1 port map( A => n12015, Z => n12014);
   U13126 : BUF_X1 port map( A => n12006, Z => n12005);
   U13127 : BUF_X1 port map( A => n11997, Z => n11996);
   U13128 : BUF_X1 port map( A => n11988, Z => n11987);
   U13129 : BUF_X1 port map( A => n11979, Z => n11978);
   U13130 : BUF_X1 port map( A => n11970, Z => n11969);
   U13131 : BUF_X1 port map( A => n11961, Z => n11960);
   U13132 : BUF_X1 port map( A => n11952, Z => n11951);
   U13133 : BUF_X1 port map( A => n11943, Z => n11942);
   U13134 : BUF_X1 port map( A => n11934, Z => n11933);
   U13135 : BUF_X1 port map( A => n11925, Z => n11924);
   U13136 : BUF_X1 port map( A => n11916, Z => n11915);
   U13137 : BUF_X1 port map( A => n11907, Z => n11906);
   U13138 : BUF_X1 port map( A => n11898, Z => n11897);
   U13139 : BUF_X1 port map( A => n11872, Z => n11667);
   U13140 : BUF_X1 port map( A => n11873, Z => n11872);
   U13141 : BUF_X1 port map( A => n11028, Z => n11027);
   U13142 : BUF_X1 port map( A => n10803, Z => n10802);
   U13143 : BUF_X1 port map( A => N4249, Z => n11891);
   U13144 : OAI21_X1 port map( B1 => n7275, B2 => n7276, A => n11508, ZN => 
                           N4249);
   U13145 : BUF_X1 port map( A => n11873, Z => n11871);
   U13146 : BUF_X1 port map( A => n11873, Z => n11870);
   U13147 : BUF_X1 port map( A => n11873, Z => n11869);
   U13148 : BUF_X1 port map( A => n11873, Z => n11868);
   U13149 : BUF_X1 port map( A => n7311, Z => n10950);
   U13150 : NAND2_X1 port map( A1 => n8462, A2 => n10995, ZN => n7311);
   U13151 : BUF_X1 port map( A => n7308, Z => n10977);
   U13152 : NAND2_X1 port map( A1 => n8462, A2 => n11012, ZN => n7308);
   U13153 : BUF_X1 port map( A => n8491, Z => n10725);
   U13154 : NAND2_X1 port map( A1 => n9642, A2 => n10770, ZN => n8491);
   U13155 : BUF_X1 port map( A => n8488, Z => n10752);
   U13156 : NAND2_X1 port map( A1 => n9642, A2 => n10787, ZN => n8488);
   U13157 : BUF_X1 port map( A => n11044, Z => n11043);
   U13158 : BUF_X1 port map( A => n11062, Z => n11061);
   U13159 : BUF_X1 port map( A => n10819, Z => n10818);
   U13160 : BUF_X1 port map( A => n10837, Z => n10836);
   U13161 : BUF_X1 port map( A => n11532, Z => n11547);
   U13162 : BUF_X1 port map( A => n6246, Z => n11532);
   U13163 : BUF_X1 port map( A => n11549, Z => n11564);
   U13164 : BUF_X1 port map( A => n6245, Z => n11549);
   U13165 : BUF_X1 port map( A => n11583, Z => n11598);
   U13166 : BUF_X1 port map( A => n6243, Z => n11583);
   U13167 : BUF_X1 port map( A => n11566, Z => n11581);
   U13168 : BUF_X1 port map( A => n6244, Z => n11566);
   U13169 : BUF_X1 port map( A => n11600, Z => n11615);
   U13170 : BUF_X1 port map( A => n6237, Z => n11600);
   U13171 : BUF_X1 port map( A => n11617, Z => n11632);
   U13172 : BUF_X1 port map( A => n6236, Z => n11617);
   U13173 : BUF_X1 port map( A => n11651, Z => n11666);
   U13174 : BUF_X1 port map( A => n6234, Z => n11651);
   U13175 : BUF_X1 port map( A => n11634, Z => n11649);
   U13176 : BUF_X1 port map( A => n6235, Z => n11634);
   U13177 : BUF_X1 port map( A => n11005, Z => n11002);
   U13178 : BUF_X1 port map( A => n11005, Z => n11003);
   U13179 : BUF_X1 port map( A => n10780, Z => n10777);
   U13180 : BUF_X1 port map( A => n10780, Z => n10778);
   U13181 : BUF_X1 port map( A => n11005, Z => n11004);
   U13182 : BUF_X1 port map( A => n10780, Z => n10779);
   U13183 : BUF_X1 port map( A => n11008, Z => n10995);
   U13184 : BUF_X1 port map( A => n11009, Z => n11008);
   U13185 : BUF_X1 port map( A => n10783, Z => n10770);
   U13186 : BUF_X1 port map( A => n10784, Z => n10783);
   U13187 : BUF_X1 port map( A => n11058, Z => n11055);
   U13188 : BUF_X1 port map( A => n11058, Z => n11056);
   U13189 : BUF_X1 port map( A => n10833, Z => n10830);
   U13190 : BUF_X1 port map( A => n10833, Z => n10831);
   U13191 : BUF_X1 port map( A => n11040, Z => n11037);
   U13192 : BUF_X1 port map( A => n11040, Z => n11038);
   U13193 : BUF_X1 port map( A => n10815, Z => n10812);
   U13194 : BUF_X1 port map( A => n10815, Z => n10813);
   U13195 : BUF_X1 port map( A => n10993, Z => n10991);
   U13196 : BUF_X1 port map( A => n10993, Z => n10990);
   U13197 : BUF_X1 port map( A => n10994, Z => n10989);
   U13198 : BUF_X1 port map( A => n10994, Z => n10988);
   U13199 : BUF_X1 port map( A => n10994, Z => n10987);
   U13200 : BUF_X1 port map( A => n10768, Z => n10766);
   U13201 : BUF_X1 port map( A => n10768, Z => n10765);
   U13202 : BUF_X1 port map( A => n10769, Z => n10764);
   U13203 : BUF_X1 port map( A => n10769, Z => n10763);
   U13204 : BUF_X1 port map( A => n10769, Z => n10762);
   U13205 : BUF_X1 port map( A => n11058, Z => n11057);
   U13206 : BUF_X1 port map( A => n10833, Z => n10832);
   U13207 : BUF_X1 port map( A => n11040, Z => n11039);
   U13208 : BUF_X1 port map( A => n10815, Z => n10814);
   U13209 : BUF_X1 port map( A => n12178, Z => n12171);
   U13210 : BUF_X1 port map( A => n12178, Z => n12172);
   U13211 : BUF_X1 port map( A => n12178, Z => n12173);
   U13212 : BUF_X1 port map( A => n12177, Z => n12174);
   U13213 : BUF_X1 port map( A => n12177, Z => n12175);
   U13214 : BUF_X1 port map( A => n12186, Z => n12179);
   U13215 : BUF_X1 port map( A => n12186, Z => n12180);
   U13216 : BUF_X1 port map( A => n12186, Z => n12181);
   U13217 : BUF_X1 port map( A => n12185, Z => n12182);
   U13218 : BUF_X1 port map( A => n12185, Z => n12183);
   U13219 : BUF_X1 port map( A => n10993, Z => n10992);
   U13220 : BUF_X1 port map( A => n10768, Z => n10767);
   U13221 : BUF_X1 port map( A => n12177, Z => n12176);
   U13222 : BUF_X1 port map( A => n12185, Z => n12184);
   U13223 : NOR2_X1 port map( A1 => n6242, A2 => n6241, ZN => n8462);
   U13224 : NOR2_X1 port map( A1 => n6233, A2 => n6232, ZN => n9642);
   U13225 : NAND2_X1 port map( A1 => n6227, A2 => n6228, ZN => n7275);
   U13226 : NOR4_X1 port map( A1 => n7290, A2 => n7291, A3 => n7292, A4 => 
                           n7293, ZN => n7289);
   U13227 : AOI221_X1 port map( B1 => n10880, B2 => n10159, C1 => n10872, C2 =>
                           n9711, A => n7324, ZN => n7287);
   U13228 : AOI221_X1 port map( B1 => n10923, B2 => n10160, C1 => n10915, C2 =>
                           n9712, A => n7318, ZN => n7288);
   U13229 : NOR4_X1 port map( A1 => n7330, A2 => n7331, A3 => n7332, A4 => 
                           n7333, ZN => n7329);
   U13230 : AOI221_X1 port map( B1 => n10880, B2 => n10161, C1 => n10872, C2 =>
                           n9713, A => n7344, ZN => n7327);
   U13231 : AOI221_X1 port map( B1 => n10923, B2 => n10162, C1 => n10915, C2 =>
                           n9714, A => n7343, ZN => n7328);
   U13232 : NOR4_X1 port map( A1 => n7348, A2 => n7349, A3 => n7350, A4 => 
                           n7351, ZN => n7347);
   U13233 : AOI221_X1 port map( B1 => n10880, B2 => n10163, C1 => n10872, C2 =>
                           n9715, A => n7362, ZN => n7345);
   U13234 : AOI221_X1 port map( B1 => n10923, B2 => n10164, C1 => n10915, C2 =>
                           n9716, A => n7361, ZN => n7346);
   U13235 : NOR4_X1 port map( A1 => n7366, A2 => n7367, A3 => n7368, A4 => 
                           n7369, ZN => n7365);
   U13236 : AOI221_X1 port map( B1 => n10880, B2 => n10165, C1 => n10872, C2 =>
                           n9717, A => n7380, ZN => n7363);
   U13237 : AOI221_X1 port map( B1 => n10923, B2 => n10166, C1 => n10915, C2 =>
                           n9718, A => n7379, ZN => n7364);
   U13238 : NOR4_X1 port map( A1 => n7384, A2 => n7385, A3 => n7386, A4 => 
                           n7387, ZN => n7383);
   U13239 : AOI221_X1 port map( B1 => n10879, B2 => n10167, C1 => n10871, C2 =>
                           n9719, A => n7398, ZN => n7381);
   U13240 : AOI221_X1 port map( B1 => n10922, B2 => n10168, C1 => n10914, C2 =>
                           n9720, A => n7397, ZN => n7382);
   U13241 : NOR4_X1 port map( A1 => n7402, A2 => n7403, A3 => n7404, A4 => 
                           n7405, ZN => n7401);
   U13242 : AOI221_X1 port map( B1 => n10879, B2 => n10169, C1 => n10871, C2 =>
                           n9721, A => n7416, ZN => n7399);
   U13243 : AOI221_X1 port map( B1 => n10922, B2 => n10170, C1 => n10914, C2 =>
                           n9722, A => n7415, ZN => n7400);
   U13244 : NOR4_X1 port map( A1 => n7420, A2 => n7421, A3 => n7422, A4 => 
                           n7423, ZN => n7419);
   U13245 : AOI221_X1 port map( B1 => n10879, B2 => n10171, C1 => n10871, C2 =>
                           n9723, A => n7434, ZN => n7417);
   U13246 : AOI221_X1 port map( B1 => n10922, B2 => n10172, C1 => n10914, C2 =>
                           n9724, A => n7433, ZN => n7418);
   U13247 : NOR4_X1 port map( A1 => n7438, A2 => n7439, A3 => n7440, A4 => 
                           n7441, ZN => n7437);
   U13248 : AOI221_X1 port map( B1 => n10879, B2 => n10173, C1 => n10871, C2 =>
                           n9725, A => n7452, ZN => n7435);
   U13249 : AOI221_X1 port map( B1 => n10922, B2 => n10174, C1 => n10914, C2 =>
                           n9726, A => n7451, ZN => n7436);
   U13250 : NOR4_X1 port map( A1 => n7456, A2 => n7457, A3 => n7458, A4 => 
                           n7459, ZN => n7455);
   U13251 : AOI221_X1 port map( B1 => n10879, B2 => n10175, C1 => n10871, C2 =>
                           n9727, A => n7470, ZN => n7453);
   U13252 : AOI221_X1 port map( B1 => n10922, B2 => n10176, C1 => n10914, C2 =>
                           n9728, A => n7469, ZN => n7454);
   U13253 : NOR4_X1 port map( A1 => n7474, A2 => n7475, A3 => n7476, A4 => 
                           n7477, ZN => n7473);
   U13254 : AOI221_X1 port map( B1 => n10879, B2 => n10177, C1 => n10871, C2 =>
                           n9729, A => n7488, ZN => n7471);
   U13255 : AOI221_X1 port map( B1 => n10922, B2 => n10178, C1 => n10914, C2 =>
                           n9730, A => n7487, ZN => n7472);
   U13256 : NOR4_X1 port map( A1 => n7492, A2 => n7493, A3 => n7494, A4 => 
                           n7495, ZN => n7491);
   U13257 : AOI221_X1 port map( B1 => n10879, B2 => n10179, C1 => n10871, C2 =>
                           n9731, A => n7506, ZN => n7489);
   U13258 : AOI221_X1 port map( B1 => n10922, B2 => n10180, C1 => n10914, C2 =>
                           n9732, A => n7505, ZN => n7490);
   U13259 : NOR4_X1 port map( A1 => n7510, A2 => n7511, A3 => n7512, A4 => 
                           n7513, ZN => n7509);
   U13260 : AOI221_X1 port map( B1 => n10879, B2 => n10181, C1 => n10871, C2 =>
                           n9733, A => n7524, ZN => n7507);
   U13261 : AOI221_X1 port map( B1 => n10922, B2 => n10182, C1 => n10914, C2 =>
                           n9734, A => n7523, ZN => n7508);
   U13262 : NOR4_X1 port map( A1 => n7528, A2 => n7529, A3 => n7530, A4 => 
                           n7531, ZN => n7527);
   U13263 : AOI221_X1 port map( B1 => n10879, B2 => n10183, C1 => n10871, C2 =>
                           n9735, A => n7542, ZN => n7525);
   U13264 : AOI221_X1 port map( B1 => n10922, B2 => n10184, C1 => n10914, C2 =>
                           n9736, A => n7541, ZN => n7526);
   U13265 : NOR4_X1 port map( A1 => n7546, A2 => n7547, A3 => n7548, A4 => 
                           n7549, ZN => n7545);
   U13266 : AOI221_X1 port map( B1 => n10879, B2 => n10185, C1 => n10871, C2 =>
                           n9737, A => n7560, ZN => n7543);
   U13267 : AOI221_X1 port map( B1 => n10922, B2 => n10186, C1 => n10914, C2 =>
                           n9738, A => n7559, ZN => n7544);
   U13268 : NOR4_X1 port map( A1 => n7564, A2 => n7565, A3 => n7566, A4 => 
                           n7567, ZN => n7563);
   U13269 : AOI221_X1 port map( B1 => n10879, B2 => n10187, C1 => n10871, C2 =>
                           n9739, A => n7578, ZN => n7561);
   U13270 : AOI221_X1 port map( B1 => n10922, B2 => n10188, C1 => n10914, C2 =>
                           n9740, A => n7577, ZN => n7562);
   U13271 : NOR4_X1 port map( A1 => n7582, A2 => n7583, A3 => n7584, A4 => 
                           n7585, ZN => n7581);
   U13272 : AOI221_X1 port map( B1 => n10879, B2 => n10189, C1 => n10871, C2 =>
                           n9741, A => n7596, ZN => n7579);
   U13273 : AOI221_X1 port map( B1 => n10922, B2 => n10190, C1 => n10914, C2 =>
                           n9742, A => n7595, ZN => n7580);
   U13274 : NOR4_X1 port map( A1 => n7600, A2 => n7601, A3 => n7602, A4 => 
                           n7603, ZN => n7599);
   U13275 : AOI221_X1 port map( B1 => n10878, B2 => n10191, C1 => n10870, C2 =>
                           n9743, A => n7614, ZN => n7597);
   U13276 : AOI221_X1 port map( B1 => n10921, B2 => n10192, C1 => n10913, C2 =>
                           n9744, A => n7613, ZN => n7598);
   U13277 : NOR4_X1 port map( A1 => n7618, A2 => n7619, A3 => n7620, A4 => 
                           n7621, ZN => n7617);
   U13278 : AOI221_X1 port map( B1 => n10878, B2 => n10193, C1 => n10870, C2 =>
                           n9745, A => n7632, ZN => n7615);
   U13279 : AOI221_X1 port map( B1 => n10921, B2 => n10194, C1 => n10913, C2 =>
                           n9746, A => n7631, ZN => n7616);
   U13280 : NOR4_X1 port map( A1 => n7636, A2 => n7637, A3 => n7638, A4 => 
                           n7639, ZN => n7635);
   U13281 : AOI221_X1 port map( B1 => n10878, B2 => n10195, C1 => n10870, C2 =>
                           n9747, A => n7650, ZN => n7633);
   U13282 : AOI221_X1 port map( B1 => n10921, B2 => n10196, C1 => n10913, C2 =>
                           n9748, A => n7649, ZN => n7634);
   U13283 : NOR4_X1 port map( A1 => n7654, A2 => n7655, A3 => n7656, A4 => 
                           n7657, ZN => n7653);
   U13284 : AOI221_X1 port map( B1 => n10878, B2 => n10197, C1 => n10870, C2 =>
                           n9749, A => n7668, ZN => n7651);
   U13285 : AOI221_X1 port map( B1 => n10921, B2 => n10198, C1 => n10913, C2 =>
                           n9750, A => n7667, ZN => n7652);
   U13286 : NOR4_X1 port map( A1 => n7672, A2 => n7673, A3 => n7674, A4 => 
                           n7675, ZN => n7671);
   U13287 : AOI221_X1 port map( B1 => n10878, B2 => n10199, C1 => n10870, C2 =>
                           n9751, A => n7686, ZN => n7669);
   U13288 : AOI221_X1 port map( B1 => n10921, B2 => n10200, C1 => n10913, C2 =>
                           n9752, A => n7685, ZN => n7670);
   U13289 : NOR4_X1 port map( A1 => n7690, A2 => n7691, A3 => n7692, A4 => 
                           n7693, ZN => n7689);
   U13290 : AOI221_X1 port map( B1 => n10878, B2 => n10201, C1 => n10870, C2 =>
                           n9753, A => n7704, ZN => n7687);
   U13291 : AOI221_X1 port map( B1 => n10921, B2 => n10202, C1 => n10913, C2 =>
                           n9754, A => n7703, ZN => n7688);
   U13292 : NOR4_X1 port map( A1 => n7708, A2 => n7709, A3 => n7710, A4 => 
                           n7711, ZN => n7707);
   U13293 : AOI221_X1 port map( B1 => n10878, B2 => n10203, C1 => n10870, C2 =>
                           n9755, A => n7722, ZN => n7705);
   U13294 : AOI221_X1 port map( B1 => n10921, B2 => n10204, C1 => n10913, C2 =>
                           n9756, A => n7721, ZN => n7706);
   U13295 : NOR4_X1 port map( A1 => n7726, A2 => n7727, A3 => n7728, A4 => 
                           n7729, ZN => n7725);
   U13296 : AOI221_X1 port map( B1 => n10878, B2 => n10205, C1 => n10870, C2 =>
                           n9757, A => n7740, ZN => n7723);
   U13297 : AOI221_X1 port map( B1 => n10921, B2 => n10206, C1 => n10913, C2 =>
                           n9758, A => n7739, ZN => n7724);
   U13298 : NOR4_X1 port map( A1 => n7744, A2 => n7745, A3 => n7746, A4 => 
                           n7747, ZN => n7743);
   U13299 : AOI221_X1 port map( B1 => n10878, B2 => n10207, C1 => n10870, C2 =>
                           n9759, A => n7758, ZN => n7741);
   U13300 : AOI221_X1 port map( B1 => n10921, B2 => n10208, C1 => n10913, C2 =>
                           n9760, A => n7757, ZN => n7742);
   U13301 : NOR4_X1 port map( A1 => n7762, A2 => n7763, A3 => n7764, A4 => 
                           n7765, ZN => n7761);
   U13302 : AOI221_X1 port map( B1 => n10878, B2 => n10209, C1 => n10870, C2 =>
                           n9761, A => n7776, ZN => n7759);
   U13303 : AOI221_X1 port map( B1 => n10921, B2 => n10210, C1 => n10913, C2 =>
                           n9762, A => n7775, ZN => n7760);
   U13304 : NOR4_X1 port map( A1 => n7780, A2 => n7781, A3 => n7782, A4 => 
                           n7783, ZN => n7779);
   U13305 : AOI221_X1 port map( B1 => n10878, B2 => n10211, C1 => n10870, C2 =>
                           n9763, A => n7794, ZN => n7777);
   U13306 : AOI221_X1 port map( B1 => n10921, B2 => n10212, C1 => n10913, C2 =>
                           n9764, A => n7793, ZN => n7778);
   U13307 : NOR4_X1 port map( A1 => n7798, A2 => n7799, A3 => n7800, A4 => 
                           n7801, ZN => n7797);
   U13308 : AOI221_X1 port map( B1 => n10878, B2 => n10213, C1 => n10870, C2 =>
                           n9765, A => n7812, ZN => n7795);
   U13309 : AOI221_X1 port map( B1 => n10921, B2 => n10214, C1 => n10913, C2 =>
                           n9766, A => n7811, ZN => n7796);
   U13310 : NOR4_X1 port map( A1 => n7816, A2 => n7817, A3 => n7818, A4 => 
                           n7819, ZN => n7815);
   U13311 : AOI221_X1 port map( B1 => n10877, B2 => n10215, C1 => n10869, C2 =>
                           n9767, A => n7830, ZN => n7813);
   U13312 : AOI221_X1 port map( B1 => n10920, B2 => n10216, C1 => n10912, C2 =>
                           n9768, A => n7829, ZN => n7814);
   U13313 : NOR4_X1 port map( A1 => n7834, A2 => n7835, A3 => n7836, A4 => 
                           n7837, ZN => n7833);
   U13314 : AOI221_X1 port map( B1 => n10877, B2 => n10217, C1 => n10869, C2 =>
                           n9769, A => n7848, ZN => n7831);
   U13315 : AOI221_X1 port map( B1 => n10920, B2 => n10218, C1 => n10912, C2 =>
                           n9770, A => n7847, ZN => n7832);
   U13316 : NOR4_X1 port map( A1 => n7852, A2 => n7853, A3 => n7854, A4 => 
                           n7855, ZN => n7851);
   U13317 : AOI221_X1 port map( B1 => n10877, B2 => n10219, C1 => n10869, C2 =>
                           n9771, A => n7866, ZN => n7849);
   U13318 : AOI221_X1 port map( B1 => n10920, B2 => n10220, C1 => n10912, C2 =>
                           n9772, A => n7865, ZN => n7850);
   U13319 : NOR4_X1 port map( A1 => n7870, A2 => n7871, A3 => n7872, A4 => 
                           n7873, ZN => n7869);
   U13320 : AOI221_X1 port map( B1 => n10877, B2 => n10221, C1 => n10869, C2 =>
                           n9773, A => n7884, ZN => n7867);
   U13321 : AOI221_X1 port map( B1 => n10920, B2 => n10222, C1 => n10912, C2 =>
                           n9774, A => n7883, ZN => n7868);
   U13322 : NOR4_X1 port map( A1 => n7888, A2 => n7889, A3 => n7890, A4 => 
                           n7891, ZN => n7887);
   U13323 : AOI221_X1 port map( B1 => n10877, B2 => n10223, C1 => n10869, C2 =>
                           n9775, A => n7902, ZN => n7885);
   U13324 : AOI221_X1 port map( B1 => n10920, B2 => n10224, C1 => n10912, C2 =>
                           n9776, A => n7901, ZN => n7886);
   U13325 : NOR4_X1 port map( A1 => n7906, A2 => n7907, A3 => n7908, A4 => 
                           n7909, ZN => n7905);
   U13326 : AOI221_X1 port map( B1 => n10877, B2 => n10225, C1 => n10869, C2 =>
                           n9777, A => n7920, ZN => n7903);
   U13327 : AOI221_X1 port map( B1 => n10920, B2 => n10226, C1 => n10912, C2 =>
                           n9778, A => n7919, ZN => n7904);
   U13328 : NOR4_X1 port map( A1 => n7924, A2 => n7925, A3 => n7926, A4 => 
                           n7927, ZN => n7923);
   U13329 : AOI221_X1 port map( B1 => n10877, B2 => n10227, C1 => n10869, C2 =>
                           n9779, A => n7938, ZN => n7921);
   U13330 : AOI221_X1 port map( B1 => n10920, B2 => n10228, C1 => n10912, C2 =>
                           n9780, A => n7937, ZN => n7922);
   U13331 : NOR4_X1 port map( A1 => n7942, A2 => n7943, A3 => n7944, A4 => 
                           n7945, ZN => n7941);
   U13332 : AOI221_X1 port map( B1 => n10877, B2 => n10229, C1 => n10869, C2 =>
                           n9781, A => n7956, ZN => n7939);
   U13333 : AOI221_X1 port map( B1 => n10920, B2 => n10230, C1 => n10912, C2 =>
                           n9782, A => n7955, ZN => n7940);
   U13334 : NOR4_X1 port map( A1 => n7960, A2 => n7961, A3 => n7962, A4 => 
                           n7963, ZN => n7959);
   U13335 : AOI221_X1 port map( B1 => n10877, B2 => n10231, C1 => n10869, C2 =>
                           n9783, A => n7974, ZN => n7957);
   U13336 : AOI221_X1 port map( B1 => n10920, B2 => n10232, C1 => n10912, C2 =>
                           n9784, A => n7973, ZN => n7958);
   U13337 : NOR4_X1 port map( A1 => n7978, A2 => n7979, A3 => n7980, A4 => 
                           n7981, ZN => n7977);
   U13338 : AOI221_X1 port map( B1 => n10877, B2 => n10233, C1 => n10869, C2 =>
                           n9785, A => n7992, ZN => n7975);
   U13339 : AOI221_X1 port map( B1 => n10920, B2 => n10234, C1 => n10912, C2 =>
                           n9786, A => n7991, ZN => n7976);
   U13340 : NOR4_X1 port map( A1 => n7996, A2 => n7997, A3 => n7998, A4 => 
                           n7999, ZN => n7995);
   U13341 : AOI221_X1 port map( B1 => n10877, B2 => n10235, C1 => n10869, C2 =>
                           n9787, A => n8010, ZN => n7993);
   U13342 : AOI221_X1 port map( B1 => n10920, B2 => n10236, C1 => n10912, C2 =>
                           n9788, A => n8009, ZN => n7994);
   U13343 : NOR4_X1 port map( A1 => n8014, A2 => n8015, A3 => n8016, A4 => 
                           n8017, ZN => n8013);
   U13344 : AOI221_X1 port map( B1 => n10877, B2 => n10237, C1 => n10869, C2 =>
                           n9789, A => n8028, ZN => n8011);
   U13345 : AOI221_X1 port map( B1 => n10920, B2 => n10238, C1 => n10912, C2 =>
                           n9790, A => n8027, ZN => n8012);
   U13346 : NOR4_X1 port map( A1 => n8032, A2 => n8033, A3 => n8034, A4 => 
                           n8035, ZN => n8031);
   U13347 : AOI221_X1 port map( B1 => n10876, B2 => n10239, C1 => n10868, C2 =>
                           n9791, A => n8046, ZN => n8029);
   U13348 : AOI221_X1 port map( B1 => n10919, B2 => n10240, C1 => n10911, C2 =>
                           n9792, A => n8045, ZN => n8030);
   U13349 : NOR4_X1 port map( A1 => n8050, A2 => n8051, A3 => n8052, A4 => 
                           n8053, ZN => n8049);
   U13350 : AOI221_X1 port map( B1 => n10876, B2 => n10241, C1 => n10868, C2 =>
                           n9793, A => n8064, ZN => n8047);
   U13351 : AOI221_X1 port map( B1 => n10919, B2 => n10242, C1 => n10911, C2 =>
                           n9794, A => n8063, ZN => n8048);
   U13352 : NOR4_X1 port map( A1 => n8068, A2 => n8069, A3 => n8070, A4 => 
                           n8071, ZN => n8067);
   U13353 : AOI221_X1 port map( B1 => n10876, B2 => n10243, C1 => n10868, C2 =>
                           n9795, A => n8082, ZN => n8065);
   U13354 : AOI221_X1 port map( B1 => n10919, B2 => n10244, C1 => n10911, C2 =>
                           n9796, A => n8081, ZN => n8066);
   U13355 : NOR4_X1 port map( A1 => n8086, A2 => n8087, A3 => n8088, A4 => 
                           n8089, ZN => n8085);
   U13356 : AOI221_X1 port map( B1 => n10876, B2 => n10245, C1 => n10868, C2 =>
                           n9797, A => n8100, ZN => n8083);
   U13357 : AOI221_X1 port map( B1 => n10919, B2 => n10246, C1 => n10911, C2 =>
                           n9798, A => n8099, ZN => n8084);
   U13358 : NOR4_X1 port map( A1 => n8104, A2 => n8105, A3 => n8106, A4 => 
                           n8107, ZN => n8103);
   U13359 : AOI221_X1 port map( B1 => n10876, B2 => n10247, C1 => n10868, C2 =>
                           n9799, A => n8118, ZN => n8101);
   U13360 : AOI221_X1 port map( B1 => n10919, B2 => n10248, C1 => n10911, C2 =>
                           n9800, A => n8117, ZN => n8102);
   U13361 : NOR4_X1 port map( A1 => n8122, A2 => n8123, A3 => n8124, A4 => 
                           n8125, ZN => n8121);
   U13362 : AOI221_X1 port map( B1 => n10876, B2 => n10249, C1 => n10868, C2 =>
                           n9801, A => n8136, ZN => n8119);
   U13363 : AOI221_X1 port map( B1 => n10919, B2 => n10250, C1 => n10911, C2 =>
                           n9802, A => n8135, ZN => n8120);
   U13364 : NOR4_X1 port map( A1 => n8140, A2 => n8141, A3 => n8142, A4 => 
                           n8143, ZN => n8139);
   U13365 : AOI221_X1 port map( B1 => n10876, B2 => n10251, C1 => n10868, C2 =>
                           n9803, A => n8154, ZN => n8137);
   U13366 : AOI221_X1 port map( B1 => n10919, B2 => n10252, C1 => n10911, C2 =>
                           n9804, A => n8153, ZN => n8138);
   U13367 : NOR4_X1 port map( A1 => n8158, A2 => n8159, A3 => n8160, A4 => 
                           n8161, ZN => n8157);
   U13368 : AOI221_X1 port map( B1 => n10876, B2 => n10253, C1 => n10868, C2 =>
                           n9805, A => n8172, ZN => n8155);
   U13369 : AOI221_X1 port map( B1 => n10919, B2 => n10254, C1 => n10911, C2 =>
                           n9806, A => n8171, ZN => n8156);
   U13370 : NOR4_X1 port map( A1 => n8176, A2 => n8177, A3 => n8178, A4 => 
                           n8179, ZN => n8175);
   U13371 : AOI221_X1 port map( B1 => n10876, B2 => n10255, C1 => n10868, C2 =>
                           n9807, A => n8190, ZN => n8173);
   U13372 : AOI221_X1 port map( B1 => n10919, B2 => n10256, C1 => n10911, C2 =>
                           n9808, A => n8189, ZN => n8174);
   U13373 : NOR4_X1 port map( A1 => n8194, A2 => n8195, A3 => n8196, A4 => 
                           n8197, ZN => n8193);
   U13374 : AOI221_X1 port map( B1 => n10876, B2 => n10257, C1 => n10868, C2 =>
                           n9809, A => n8208, ZN => n8191);
   U13375 : AOI221_X1 port map( B1 => n10919, B2 => n10258, C1 => n10911, C2 =>
                           n9810, A => n8207, ZN => n8192);
   U13376 : NOR4_X1 port map( A1 => n8212, A2 => n8213, A3 => n8214, A4 => 
                           n8215, ZN => n8211);
   U13377 : AOI221_X1 port map( B1 => n10876, B2 => n10259, C1 => n10868, C2 =>
                           n9811, A => n8226, ZN => n8209);
   U13378 : AOI221_X1 port map( B1 => n10919, B2 => n10260, C1 => n10911, C2 =>
                           n9812, A => n8225, ZN => n8210);
   U13379 : NOR4_X1 port map( A1 => n8230, A2 => n8231, A3 => n8232, A4 => 
                           n8233, ZN => n8229);
   U13380 : AOI221_X1 port map( B1 => n10876, B2 => n10261, C1 => n10868, C2 =>
                           n9813, A => n8244, ZN => n8227);
   U13381 : AOI221_X1 port map( B1 => n10919, B2 => n10262, C1 => n10911, C2 =>
                           n9814, A => n8243, ZN => n8228);
   U13382 : NOR4_X1 port map( A1 => n8248, A2 => n8249, A3 => n8250, A4 => 
                           n8251, ZN => n8247);
   U13383 : AOI221_X1 port map( B1 => n10875, B2 => n10263, C1 => n10867, C2 =>
                           n9815, A => n8262, ZN => n8245);
   U13384 : AOI221_X1 port map( B1 => n10918, B2 => n10264, C1 => n10910, C2 =>
                           n9816, A => n8261, ZN => n8246);
   U13385 : NOR4_X1 port map( A1 => n8266, A2 => n8267, A3 => n8268, A4 => 
                           n8269, ZN => n8265);
   U13386 : AOI221_X1 port map( B1 => n10875, B2 => n10265, C1 => n10867, C2 =>
                           n9817, A => n8280, ZN => n8263);
   U13387 : AOI221_X1 port map( B1 => n10918, B2 => n10266, C1 => n10910, C2 =>
                           n9818, A => n8279, ZN => n8264);
   U13388 : NOR4_X1 port map( A1 => n8284, A2 => n8285, A3 => n8286, A4 => 
                           n8287, ZN => n8283);
   U13389 : AOI221_X1 port map( B1 => n10875, B2 => n10267, C1 => n10867, C2 =>
                           n9819, A => n8298, ZN => n8281);
   U13390 : AOI221_X1 port map( B1 => n10918, B2 => n10268, C1 => n10910, C2 =>
                           n9820, A => n8297, ZN => n8282);
   U13391 : NOR4_X1 port map( A1 => n8302, A2 => n8303, A3 => n8304, A4 => 
                           n8305, ZN => n8301);
   U13392 : AOI221_X1 port map( B1 => n10875, B2 => n10269, C1 => n10867, C2 =>
                           n9821, A => n8316, ZN => n8299);
   U13393 : AOI221_X1 port map( B1 => n10918, B2 => n10270, C1 => n10910, C2 =>
                           n9822, A => n8315, ZN => n8300);
   U13394 : NOR4_X1 port map( A1 => n8320, A2 => n8321, A3 => n8322, A4 => 
                           n8323, ZN => n8319);
   U13395 : AOI221_X1 port map( B1 => n10875, B2 => n10271, C1 => n10867, C2 =>
                           n9823, A => n8334, ZN => n8317);
   U13396 : AOI221_X1 port map( B1 => n10918, B2 => n10272, C1 => n10910, C2 =>
                           n9824, A => n8333, ZN => n8318);
   U13397 : NOR4_X1 port map( A1 => n8338, A2 => n8339, A3 => n8340, A4 => 
                           n8341, ZN => n8337);
   U13398 : AOI221_X1 port map( B1 => n10875, B2 => n10273, C1 => n10867, C2 =>
                           n9825, A => n8352, ZN => n8335);
   U13399 : AOI221_X1 port map( B1 => n10918, B2 => n10274, C1 => n10910, C2 =>
                           n9826, A => n8351, ZN => n8336);
   U13400 : NOR4_X1 port map( A1 => n8356, A2 => n8357, A3 => n8358, A4 => 
                           n8359, ZN => n8355);
   U13401 : AOI221_X1 port map( B1 => n10875, B2 => n10275, C1 => n10867, C2 =>
                           n9827, A => n8370, ZN => n8353);
   U13402 : AOI221_X1 port map( B1 => n10918, B2 => n10276, C1 => n10910, C2 =>
                           n9828, A => n8369, ZN => n8354);
   U13403 : NOR4_X1 port map( A1 => n8374, A2 => n8375, A3 => n8376, A4 => 
                           n8377, ZN => n8373);
   U13404 : AOI221_X1 port map( B1 => n10875, B2 => n10277, C1 => n10867, C2 =>
                           n9829, A => n8388, ZN => n8371);
   U13405 : AOI221_X1 port map( B1 => n10918, B2 => n10278, C1 => n10910, C2 =>
                           n9830, A => n8387, ZN => n8372);
   U13406 : NOR4_X1 port map( A1 => n8392, A2 => n8393, A3 => n8394, A4 => 
                           n8395, ZN => n8391);
   U13407 : AOI221_X1 port map( B1 => n10875, B2 => n10279, C1 => n10867, C2 =>
                           n9831, A => n8406, ZN => n8389);
   U13408 : AOI221_X1 port map( B1 => n10918, B2 => n10280, C1 => n10910, C2 =>
                           n9832, A => n8405, ZN => n8390);
   U13409 : NOR4_X1 port map( A1 => n8410, A2 => n8411, A3 => n8412, A4 => 
                           n8413, ZN => n8409);
   U13410 : AOI221_X1 port map( B1 => n10875, B2 => n10281, C1 => n10867, C2 =>
                           n9833, A => n8424, ZN => n8407);
   U13411 : AOI221_X1 port map( B1 => n10918, B2 => n10282, C1 => n10910, C2 =>
                           n9834, A => n8423, ZN => n8408);
   U13412 : NOR4_X1 port map( A1 => n8428, A2 => n8429, A3 => n8430, A4 => 
                           n8431, ZN => n8427);
   U13413 : AOI221_X1 port map( B1 => n10875, B2 => n10283, C1 => n10867, C2 =>
                           n9835, A => n8442, ZN => n8425);
   U13414 : AOI221_X1 port map( B1 => n10918, B2 => n10284, C1 => n10910, C2 =>
                           n9836, A => n8441, ZN => n8426);
   U13415 : NOR4_X1 port map( A1 => n8446, A2 => n8447, A3 => n8448, A4 => 
                           n8449, ZN => n8445);
   U13416 : AOI221_X1 port map( B1 => n10875, B2 => n10285, C1 => n10867, C2 =>
                           n9837, A => n8466, ZN => n8443);
   U13417 : AOI221_X1 port map( B1 => n10918, B2 => n10286, C1 => n10910, C2 =>
                           n9838, A => n8464, ZN => n8444);
   U13418 : NOR4_X1 port map( A1 => n8470, A2 => n8471, A3 => n8472, A4 => 
                           n8473, ZN => n8469);
   U13419 : AOI221_X1 port map( B1 => n10655, B2 => n10159, C1 => n10647, C2 =>
                           n9711, A => n8504, ZN => n8467);
   U13420 : AOI221_X1 port map( B1 => n10698, B2 => n10160, C1 => n10690, C2 =>
                           n9712, A => n8498, ZN => n8468);
   U13421 : NOR4_X1 port map( A1 => n8510, A2 => n8511, A3 => n8512, A4 => 
                           n8513, ZN => n8509);
   U13422 : AOI221_X1 port map( B1 => n10655, B2 => n10161, C1 => n10647, C2 =>
                           n9713, A => n8524, ZN => n8507);
   U13423 : AOI221_X1 port map( B1 => n10698, B2 => n10162, C1 => n10690, C2 =>
                           n9714, A => n8523, ZN => n8508);
   U13424 : NOR4_X1 port map( A1 => n8528, A2 => n8529, A3 => n8530, A4 => 
                           n8531, ZN => n8527);
   U13425 : AOI221_X1 port map( B1 => n10655, B2 => n10163, C1 => n10647, C2 =>
                           n9715, A => n8542, ZN => n8525);
   U13426 : AOI221_X1 port map( B1 => n10698, B2 => n10164, C1 => n10690, C2 =>
                           n9716, A => n8541, ZN => n8526);
   U13427 : NOR4_X1 port map( A1 => n8546, A2 => n8547, A3 => n8548, A4 => 
                           n8549, ZN => n8545);
   U13428 : AOI221_X1 port map( B1 => n10655, B2 => n10165, C1 => n10647, C2 =>
                           n9717, A => n8560, ZN => n8543);
   U13429 : AOI221_X1 port map( B1 => n10698, B2 => n10166, C1 => n10690, C2 =>
                           n9718, A => n8559, ZN => n8544);
   U13430 : NOR4_X1 port map( A1 => n8564, A2 => n8565, A3 => n8566, A4 => 
                           n8567, ZN => n8563);
   U13431 : AOI221_X1 port map( B1 => n10654, B2 => n10167, C1 => n10646, C2 =>
                           n9719, A => n8578, ZN => n8561);
   U13432 : AOI221_X1 port map( B1 => n10697, B2 => n10168, C1 => n10689, C2 =>
                           n9720, A => n8577, ZN => n8562);
   U13433 : NOR4_X1 port map( A1 => n8582, A2 => n8583, A3 => n8584, A4 => 
                           n8585, ZN => n8581);
   U13434 : AOI221_X1 port map( B1 => n10654, B2 => n10169, C1 => n10646, C2 =>
                           n9721, A => n8596, ZN => n8579);
   U13435 : AOI221_X1 port map( B1 => n10697, B2 => n10170, C1 => n10689, C2 =>
                           n9722, A => n8595, ZN => n8580);
   U13436 : NOR4_X1 port map( A1 => n8600, A2 => n8601, A3 => n8602, A4 => 
                           n8603, ZN => n8599);
   U13437 : AOI221_X1 port map( B1 => n10654, B2 => n10171, C1 => n10646, C2 =>
                           n9723, A => n8614, ZN => n8597);
   U13438 : AOI221_X1 port map( B1 => n10697, B2 => n10172, C1 => n10689, C2 =>
                           n9724, A => n8613, ZN => n8598);
   U13439 : NOR4_X1 port map( A1 => n8618, A2 => n8619, A3 => n8620, A4 => 
                           n8621, ZN => n8617);
   U13440 : AOI221_X1 port map( B1 => n10654, B2 => n10173, C1 => n10646, C2 =>
                           n9725, A => n8632, ZN => n8615);
   U13441 : AOI221_X1 port map( B1 => n10697, B2 => n10174, C1 => n10689, C2 =>
                           n9726, A => n8631, ZN => n8616);
   U13442 : NOR4_X1 port map( A1 => n8636, A2 => n8637, A3 => n8638, A4 => 
                           n8639, ZN => n8635);
   U13443 : AOI221_X1 port map( B1 => n10654, B2 => n10175, C1 => n10646, C2 =>
                           n9727, A => n8650, ZN => n8633);
   U13444 : AOI221_X1 port map( B1 => n10697, B2 => n10176, C1 => n10689, C2 =>
                           n9728, A => n8649, ZN => n8634);
   U13445 : NOR4_X1 port map( A1 => n8654, A2 => n8655, A3 => n8656, A4 => 
                           n8657, ZN => n8653);
   U13446 : AOI221_X1 port map( B1 => n10654, B2 => n10177, C1 => n10646, C2 =>
                           n9729, A => n8668, ZN => n8651);
   U13447 : AOI221_X1 port map( B1 => n10697, B2 => n10178, C1 => n10689, C2 =>
                           n9730, A => n8667, ZN => n8652);
   U13448 : NOR4_X1 port map( A1 => n8672, A2 => n8673, A3 => n8674, A4 => 
                           n8675, ZN => n8671);
   U13449 : AOI221_X1 port map( B1 => n10654, B2 => n10179, C1 => n10646, C2 =>
                           n9731, A => n8686, ZN => n8669);
   U13450 : AOI221_X1 port map( B1 => n10697, B2 => n10180, C1 => n10689, C2 =>
                           n9732, A => n8685, ZN => n8670);
   U13451 : NOR4_X1 port map( A1 => n8690, A2 => n8691, A3 => n8692, A4 => 
                           n8693, ZN => n8689);
   U13452 : AOI221_X1 port map( B1 => n10654, B2 => n10181, C1 => n10646, C2 =>
                           n9733, A => n8704, ZN => n8687);
   U13453 : AOI221_X1 port map( B1 => n10697, B2 => n10182, C1 => n10689, C2 =>
                           n9734, A => n8703, ZN => n8688);
   U13454 : NOR4_X1 port map( A1 => n8708, A2 => n8709, A3 => n8710, A4 => 
                           n8711, ZN => n8707);
   U13455 : AOI221_X1 port map( B1 => n10654, B2 => n10183, C1 => n10646, C2 =>
                           n9735, A => n8722, ZN => n8705);
   U13456 : AOI221_X1 port map( B1 => n10697, B2 => n10184, C1 => n10689, C2 =>
                           n9736, A => n8721, ZN => n8706);
   U13457 : NOR4_X1 port map( A1 => n8726, A2 => n8727, A3 => n8728, A4 => 
                           n8729, ZN => n8725);
   U13458 : AOI221_X1 port map( B1 => n10654, B2 => n10185, C1 => n10646, C2 =>
                           n9737, A => n8740, ZN => n8723);
   U13459 : AOI221_X1 port map( B1 => n10697, B2 => n10186, C1 => n10689, C2 =>
                           n9738, A => n8739, ZN => n8724);
   U13460 : NOR4_X1 port map( A1 => n8744, A2 => n8745, A3 => n8746, A4 => 
                           n8747, ZN => n8743);
   U13461 : AOI221_X1 port map( B1 => n10654, B2 => n10187, C1 => n10646, C2 =>
                           n9739, A => n8758, ZN => n8741);
   U13462 : AOI221_X1 port map( B1 => n10697, B2 => n10188, C1 => n10689, C2 =>
                           n9740, A => n8757, ZN => n8742);
   U13463 : NOR4_X1 port map( A1 => n8762, A2 => n8763, A3 => n8764, A4 => 
                           n8765, ZN => n8761);
   U13464 : AOI221_X1 port map( B1 => n10654, B2 => n10189, C1 => n10646, C2 =>
                           n9741, A => n8776, ZN => n8759);
   U13465 : AOI221_X1 port map( B1 => n10697, B2 => n10190, C1 => n10689, C2 =>
                           n9742, A => n8775, ZN => n8760);
   U13466 : NOR4_X1 port map( A1 => n8780, A2 => n8781, A3 => n8782, A4 => 
                           n8783, ZN => n8779);
   U13467 : AOI221_X1 port map( B1 => n10653, B2 => n10191, C1 => n10645, C2 =>
                           n9743, A => n8794, ZN => n8777);
   U13468 : AOI221_X1 port map( B1 => n10696, B2 => n10192, C1 => n10688, C2 =>
                           n9744, A => n8793, ZN => n8778);
   U13469 : NOR4_X1 port map( A1 => n8798, A2 => n8799, A3 => n8800, A4 => 
                           n8801, ZN => n8797);
   U13470 : AOI221_X1 port map( B1 => n10653, B2 => n10193, C1 => n10645, C2 =>
                           n9745, A => n8812, ZN => n8795);
   U13471 : AOI221_X1 port map( B1 => n10696, B2 => n10194, C1 => n10688, C2 =>
                           n9746, A => n8811, ZN => n8796);
   U13472 : NOR4_X1 port map( A1 => n8816, A2 => n8817, A3 => n8818, A4 => 
                           n8819, ZN => n8815);
   U13473 : AOI221_X1 port map( B1 => n10653, B2 => n10195, C1 => n10645, C2 =>
                           n9747, A => n8830, ZN => n8813);
   U13474 : AOI221_X1 port map( B1 => n10696, B2 => n10196, C1 => n10688, C2 =>
                           n9748, A => n8829, ZN => n8814);
   U13475 : NOR4_X1 port map( A1 => n8834, A2 => n8835, A3 => n8836, A4 => 
                           n8837, ZN => n8833);
   U13476 : AOI221_X1 port map( B1 => n10653, B2 => n10197, C1 => n10645, C2 =>
                           n9749, A => n8848, ZN => n8831);
   U13477 : AOI221_X1 port map( B1 => n10696, B2 => n10198, C1 => n10688, C2 =>
                           n9750, A => n8847, ZN => n8832);
   U13478 : NOR4_X1 port map( A1 => n8852, A2 => n8853, A3 => n8854, A4 => 
                           n8855, ZN => n8851);
   U13479 : AOI221_X1 port map( B1 => n10653, B2 => n10199, C1 => n10645, C2 =>
                           n9751, A => n8866, ZN => n8849);
   U13480 : AOI221_X1 port map( B1 => n10696, B2 => n10200, C1 => n10688, C2 =>
                           n9752, A => n8865, ZN => n8850);
   U13481 : NOR4_X1 port map( A1 => n8870, A2 => n8871, A3 => n8872, A4 => 
                           n8873, ZN => n8869);
   U13482 : AOI221_X1 port map( B1 => n10653, B2 => n10201, C1 => n10645, C2 =>
                           n9753, A => n8884, ZN => n8867);
   U13483 : AOI221_X1 port map( B1 => n10696, B2 => n10202, C1 => n10688, C2 =>
                           n9754, A => n8883, ZN => n8868);
   U13484 : NOR4_X1 port map( A1 => n8888, A2 => n8889, A3 => n8890, A4 => 
                           n8891, ZN => n8887);
   U13485 : AOI221_X1 port map( B1 => n10653, B2 => n10203, C1 => n10645, C2 =>
                           n9755, A => n8902, ZN => n8885);
   U13486 : AOI221_X1 port map( B1 => n10696, B2 => n10204, C1 => n10688, C2 =>
                           n9756, A => n8901, ZN => n8886);
   U13487 : NOR4_X1 port map( A1 => n8906, A2 => n8907, A3 => n8908, A4 => 
                           n8909, ZN => n8905);
   U13488 : AOI221_X1 port map( B1 => n10653, B2 => n10205, C1 => n10645, C2 =>
                           n9757, A => n8920, ZN => n8903);
   U13489 : AOI221_X1 port map( B1 => n10696, B2 => n10206, C1 => n10688, C2 =>
                           n9758, A => n8919, ZN => n8904);
   U13490 : NOR4_X1 port map( A1 => n8924, A2 => n8925, A3 => n8926, A4 => 
                           n8927, ZN => n8923);
   U13491 : AOI221_X1 port map( B1 => n10653, B2 => n10207, C1 => n10645, C2 =>
                           n9759, A => n8938, ZN => n8921);
   U13492 : AOI221_X1 port map( B1 => n10696, B2 => n10208, C1 => n10688, C2 =>
                           n9760, A => n8937, ZN => n8922);
   U13493 : NOR4_X1 port map( A1 => n8942, A2 => n8943, A3 => n8944, A4 => 
                           n8945, ZN => n8941);
   U13494 : AOI221_X1 port map( B1 => n10653, B2 => n10209, C1 => n10645, C2 =>
                           n9761, A => n8956, ZN => n8939);
   U13495 : AOI221_X1 port map( B1 => n10696, B2 => n10210, C1 => n10688, C2 =>
                           n9762, A => n8955, ZN => n8940);
   U13496 : NOR4_X1 port map( A1 => n8960, A2 => n8961, A3 => n8962, A4 => 
                           n8963, ZN => n8959);
   U13497 : AOI221_X1 port map( B1 => n10653, B2 => n10211, C1 => n10645, C2 =>
                           n9763, A => n8974, ZN => n8957);
   U13498 : AOI221_X1 port map( B1 => n10696, B2 => n10212, C1 => n10688, C2 =>
                           n9764, A => n8973, ZN => n8958);
   U13499 : NOR4_X1 port map( A1 => n8978, A2 => n8979, A3 => n8980, A4 => 
                           n8981, ZN => n8977);
   U13500 : AOI221_X1 port map( B1 => n10653, B2 => n10213, C1 => n10645, C2 =>
                           n9765, A => n8992, ZN => n8975);
   U13501 : AOI221_X1 port map( B1 => n10696, B2 => n10214, C1 => n10688, C2 =>
                           n9766, A => n8991, ZN => n8976);
   U13502 : NOR4_X1 port map( A1 => n8996, A2 => n8997, A3 => n8998, A4 => 
                           n8999, ZN => n8995);
   U13503 : AOI221_X1 port map( B1 => n10652, B2 => n10215, C1 => n10644, C2 =>
                           n9767, A => n9010, ZN => n8993);
   U13504 : AOI221_X1 port map( B1 => n10695, B2 => n10216, C1 => n10687, C2 =>
                           n9768, A => n9009, ZN => n8994);
   U13505 : NOR4_X1 port map( A1 => n9014, A2 => n9015, A3 => n9016, A4 => 
                           n9017, ZN => n9013);
   U13506 : AOI221_X1 port map( B1 => n10652, B2 => n10217, C1 => n10644, C2 =>
                           n9769, A => n9028, ZN => n9011);
   U13507 : AOI221_X1 port map( B1 => n10695, B2 => n10218, C1 => n10687, C2 =>
                           n9770, A => n9027, ZN => n9012);
   U13508 : NOR4_X1 port map( A1 => n9032, A2 => n9033, A3 => n9034, A4 => 
                           n9035, ZN => n9031);
   U13509 : AOI221_X1 port map( B1 => n10652, B2 => n10219, C1 => n10644, C2 =>
                           n9771, A => n9046, ZN => n9029);
   U13510 : AOI221_X1 port map( B1 => n10695, B2 => n10220, C1 => n10687, C2 =>
                           n9772, A => n9045, ZN => n9030);
   U13511 : NOR4_X1 port map( A1 => n9050, A2 => n9051, A3 => n9052, A4 => 
                           n9053, ZN => n9049);
   U13512 : AOI221_X1 port map( B1 => n10652, B2 => n10221, C1 => n10644, C2 =>
                           n9773, A => n9064, ZN => n9047);
   U13513 : AOI221_X1 port map( B1 => n10695, B2 => n10222, C1 => n10687, C2 =>
                           n9774, A => n9063, ZN => n9048);
   U13514 : NOR4_X1 port map( A1 => n9068, A2 => n9069, A3 => n9070, A4 => 
                           n9071, ZN => n9067);
   U13515 : AOI221_X1 port map( B1 => n10652, B2 => n10223, C1 => n10644, C2 =>
                           n9775, A => n9082, ZN => n9065);
   U13516 : AOI221_X1 port map( B1 => n10695, B2 => n10224, C1 => n10687, C2 =>
                           n9776, A => n9081, ZN => n9066);
   U13517 : NOR4_X1 port map( A1 => n9086, A2 => n9087, A3 => n9088, A4 => 
                           n9089, ZN => n9085);
   U13518 : AOI221_X1 port map( B1 => n10652, B2 => n10225, C1 => n10644, C2 =>
                           n9777, A => n9100, ZN => n9083);
   U13519 : AOI221_X1 port map( B1 => n10695, B2 => n10226, C1 => n10687, C2 =>
                           n9778, A => n9099, ZN => n9084);
   U13520 : NOR4_X1 port map( A1 => n9104, A2 => n9105, A3 => n9106, A4 => 
                           n9107, ZN => n9103);
   U13521 : AOI221_X1 port map( B1 => n10652, B2 => n10227, C1 => n10644, C2 =>
                           n9779, A => n9118, ZN => n9101);
   U13522 : AOI221_X1 port map( B1 => n10695, B2 => n10228, C1 => n10687, C2 =>
                           n9780, A => n9117, ZN => n9102);
   U13523 : NOR4_X1 port map( A1 => n9122, A2 => n9123, A3 => n9124, A4 => 
                           n9125, ZN => n9121);
   U13524 : AOI221_X1 port map( B1 => n10652, B2 => n10229, C1 => n10644, C2 =>
                           n9781, A => n9136, ZN => n9119);
   U13525 : AOI221_X1 port map( B1 => n10695, B2 => n10230, C1 => n10687, C2 =>
                           n9782, A => n9135, ZN => n9120);
   U13526 : NOR4_X1 port map( A1 => n9140, A2 => n9141, A3 => n9142, A4 => 
                           n9143, ZN => n9139);
   U13527 : AOI221_X1 port map( B1 => n10652, B2 => n10231, C1 => n10644, C2 =>
                           n9783, A => n9154, ZN => n9137);
   U13528 : AOI221_X1 port map( B1 => n10695, B2 => n10232, C1 => n10687, C2 =>
                           n9784, A => n9153, ZN => n9138);
   U13529 : NOR4_X1 port map( A1 => n9158, A2 => n9159, A3 => n9160, A4 => 
                           n9161, ZN => n9157);
   U13530 : AOI221_X1 port map( B1 => n10652, B2 => n10233, C1 => n10644, C2 =>
                           n9785, A => n9172, ZN => n9155);
   U13531 : AOI221_X1 port map( B1 => n10695, B2 => n10234, C1 => n10687, C2 =>
                           n9786, A => n9171, ZN => n9156);
   U13532 : NOR4_X1 port map( A1 => n9176, A2 => n9177, A3 => n9178, A4 => 
                           n9179, ZN => n9175);
   U13533 : AOI221_X1 port map( B1 => n10652, B2 => n10235, C1 => n10644, C2 =>
                           n9787, A => n9190, ZN => n9173);
   U13534 : AOI221_X1 port map( B1 => n10695, B2 => n10236, C1 => n10687, C2 =>
                           n9788, A => n9189, ZN => n9174);
   U13535 : NOR4_X1 port map( A1 => n9194, A2 => n9195, A3 => n9196, A4 => 
                           n9197, ZN => n9193);
   U13536 : AOI221_X1 port map( B1 => n10652, B2 => n10237, C1 => n10644, C2 =>
                           n9789, A => n9208, ZN => n9191);
   U13537 : AOI221_X1 port map( B1 => n10695, B2 => n10238, C1 => n10687, C2 =>
                           n9790, A => n9207, ZN => n9192);
   U13538 : NOR4_X1 port map( A1 => n9212, A2 => n9213, A3 => n9214, A4 => 
                           n9215, ZN => n9211);
   U13539 : AOI221_X1 port map( B1 => n10651, B2 => n10239, C1 => n10643, C2 =>
                           n9791, A => n9226, ZN => n9209);
   U13540 : AOI221_X1 port map( B1 => n10694, B2 => n10240, C1 => n10686, C2 =>
                           n9792, A => n9225, ZN => n9210);
   U13541 : NOR4_X1 port map( A1 => n9230, A2 => n9231, A3 => n9232, A4 => 
                           n9233, ZN => n9229);
   U13542 : AOI221_X1 port map( B1 => n10651, B2 => n10241, C1 => n10643, C2 =>
                           n9793, A => n9244, ZN => n9227);
   U13543 : AOI221_X1 port map( B1 => n10694, B2 => n10242, C1 => n10686, C2 =>
                           n9794, A => n9243, ZN => n9228);
   U13544 : NOR4_X1 port map( A1 => n9248, A2 => n9249, A3 => n9250, A4 => 
                           n9251, ZN => n9247);
   U13545 : AOI221_X1 port map( B1 => n10651, B2 => n10243, C1 => n10643, C2 =>
                           n9795, A => n9262, ZN => n9245);
   U13546 : AOI221_X1 port map( B1 => n10694, B2 => n10244, C1 => n10686, C2 =>
                           n9796, A => n9261, ZN => n9246);
   U13547 : NOR4_X1 port map( A1 => n9266, A2 => n9267, A3 => n9268, A4 => 
                           n9269, ZN => n9265);
   U13548 : AOI221_X1 port map( B1 => n10651, B2 => n10245, C1 => n10643, C2 =>
                           n9797, A => n9280, ZN => n9263);
   U13549 : AOI221_X1 port map( B1 => n10694, B2 => n10246, C1 => n10686, C2 =>
                           n9798, A => n9279, ZN => n9264);
   U13550 : NOR4_X1 port map( A1 => n9284, A2 => n9285, A3 => n9286, A4 => 
                           n9287, ZN => n9283);
   U13551 : AOI221_X1 port map( B1 => n10651, B2 => n10247, C1 => n10643, C2 =>
                           n9799, A => n9298, ZN => n9281);
   U13552 : AOI221_X1 port map( B1 => n10694, B2 => n10248, C1 => n10686, C2 =>
                           n9800, A => n9297, ZN => n9282);
   U13553 : NOR4_X1 port map( A1 => n9302, A2 => n9303, A3 => n9304, A4 => 
                           n9305, ZN => n9301);
   U13554 : AOI221_X1 port map( B1 => n10651, B2 => n10249, C1 => n10643, C2 =>
                           n9801, A => n9316, ZN => n9299);
   U13555 : AOI221_X1 port map( B1 => n10694, B2 => n10250, C1 => n10686, C2 =>
                           n9802, A => n9315, ZN => n9300);
   U13556 : NOR4_X1 port map( A1 => n9320, A2 => n9321, A3 => n9322, A4 => 
                           n9323, ZN => n9319);
   U13557 : AOI221_X1 port map( B1 => n10651, B2 => n10251, C1 => n10643, C2 =>
                           n9803, A => n9334, ZN => n9317);
   U13558 : AOI221_X1 port map( B1 => n10694, B2 => n10252, C1 => n10686, C2 =>
                           n9804, A => n9333, ZN => n9318);
   U13559 : NOR4_X1 port map( A1 => n9338, A2 => n9339, A3 => n9340, A4 => 
                           n9341, ZN => n9337);
   U13560 : AOI221_X1 port map( B1 => n10651, B2 => n10253, C1 => n10643, C2 =>
                           n9805, A => n9352, ZN => n9335);
   U13561 : AOI221_X1 port map( B1 => n10694, B2 => n10254, C1 => n10686, C2 =>
                           n9806, A => n9351, ZN => n9336);
   U13562 : NOR4_X1 port map( A1 => n9356, A2 => n9357, A3 => n9358, A4 => 
                           n9359, ZN => n9355);
   U13563 : AOI221_X1 port map( B1 => n10651, B2 => n10255, C1 => n10643, C2 =>
                           n9807, A => n9370, ZN => n9353);
   U13564 : AOI221_X1 port map( B1 => n10694, B2 => n10256, C1 => n10686, C2 =>
                           n9808, A => n9369, ZN => n9354);
   U13565 : NOR4_X1 port map( A1 => n9374, A2 => n9375, A3 => n9376, A4 => 
                           n9377, ZN => n9373);
   U13566 : AOI221_X1 port map( B1 => n10651, B2 => n10257, C1 => n10643, C2 =>
                           n9809, A => n9388, ZN => n9371);
   U13567 : AOI221_X1 port map( B1 => n10694, B2 => n10258, C1 => n10686, C2 =>
                           n9810, A => n9387, ZN => n9372);
   U13568 : NOR4_X1 port map( A1 => n9392, A2 => n9393, A3 => n9394, A4 => 
                           n9395, ZN => n9391);
   U13569 : AOI221_X1 port map( B1 => n10651, B2 => n10259, C1 => n10643, C2 =>
                           n9811, A => n9406, ZN => n9389);
   U13570 : AOI221_X1 port map( B1 => n10694, B2 => n10260, C1 => n10686, C2 =>
                           n9812, A => n9405, ZN => n9390);
   U13571 : NOR4_X1 port map( A1 => n9410, A2 => n9411, A3 => n9412, A4 => 
                           n9413, ZN => n9409);
   U13572 : AOI221_X1 port map( B1 => n10651, B2 => n10261, C1 => n10643, C2 =>
                           n9813, A => n9424, ZN => n9407);
   U13573 : AOI221_X1 port map( B1 => n10694, B2 => n10262, C1 => n10686, C2 =>
                           n9814, A => n9423, ZN => n9408);
   U13574 : NOR4_X1 port map( A1 => n9428, A2 => n9429, A3 => n9430, A4 => 
                           n9431, ZN => n9427);
   U13575 : AOI221_X1 port map( B1 => n10650, B2 => n10263, C1 => n10642, C2 =>
                           n9815, A => n9442, ZN => n9425);
   U13576 : AOI221_X1 port map( B1 => n10693, B2 => n10264, C1 => n10685, C2 =>
                           n9816, A => n9441, ZN => n9426);
   U13577 : NOR4_X1 port map( A1 => n9446, A2 => n9447, A3 => n9448, A4 => 
                           n9449, ZN => n9445);
   U13578 : AOI221_X1 port map( B1 => n10650, B2 => n10265, C1 => n10642, C2 =>
                           n9817, A => n9460, ZN => n9443);
   U13579 : AOI221_X1 port map( B1 => n10693, B2 => n10266, C1 => n10685, C2 =>
                           n9818, A => n9459, ZN => n9444);
   U13580 : NOR4_X1 port map( A1 => n9464, A2 => n9465, A3 => n9466, A4 => 
                           n9467, ZN => n9463);
   U13581 : AOI221_X1 port map( B1 => n10650, B2 => n10267, C1 => n10642, C2 =>
                           n9819, A => n9478, ZN => n9461);
   U13582 : AOI221_X1 port map( B1 => n10693, B2 => n10268, C1 => n10685, C2 =>
                           n9820, A => n9477, ZN => n9462);
   U13583 : NOR4_X1 port map( A1 => n9482, A2 => n9483, A3 => n9484, A4 => 
                           n9485, ZN => n9481);
   U13584 : AOI221_X1 port map( B1 => n10650, B2 => n10269, C1 => n10642, C2 =>
                           n9821, A => n9496, ZN => n9479);
   U13585 : AOI221_X1 port map( B1 => n10693, B2 => n10270, C1 => n10685, C2 =>
                           n9822, A => n9495, ZN => n9480);
   U13586 : NOR4_X1 port map( A1 => n9500, A2 => n9501, A3 => n9502, A4 => 
                           n9503, ZN => n9499);
   U13587 : AOI221_X1 port map( B1 => n10650, B2 => n10271, C1 => n10642, C2 =>
                           n9823, A => n9514, ZN => n9497);
   U13588 : AOI221_X1 port map( B1 => n10693, B2 => n10272, C1 => n10685, C2 =>
                           n9824, A => n9513, ZN => n9498);
   U13589 : NOR4_X1 port map( A1 => n9518, A2 => n9519, A3 => n9520, A4 => 
                           n9521, ZN => n9517);
   U13590 : AOI221_X1 port map( B1 => n10650, B2 => n10273, C1 => n10642, C2 =>
                           n9825, A => n9532, ZN => n9515);
   U13591 : AOI221_X1 port map( B1 => n10693, B2 => n10274, C1 => n10685, C2 =>
                           n9826, A => n9531, ZN => n9516);
   U13592 : NOR4_X1 port map( A1 => n9536, A2 => n9537, A3 => n9538, A4 => 
                           n9539, ZN => n9535);
   U13593 : AOI221_X1 port map( B1 => n10650, B2 => n10275, C1 => n10642, C2 =>
                           n9827, A => n9550, ZN => n9533);
   U13594 : AOI221_X1 port map( B1 => n10693, B2 => n10276, C1 => n10685, C2 =>
                           n9828, A => n9549, ZN => n9534);
   U13595 : NOR4_X1 port map( A1 => n9554, A2 => n9555, A3 => n9556, A4 => 
                           n9557, ZN => n9553);
   U13596 : AOI221_X1 port map( B1 => n10650, B2 => n10277, C1 => n10642, C2 =>
                           n9829, A => n9568, ZN => n9551);
   U13597 : AOI221_X1 port map( B1 => n10693, B2 => n10278, C1 => n10685, C2 =>
                           n9830, A => n9567, ZN => n9552);
   U13598 : NOR4_X1 port map( A1 => n9572, A2 => n9573, A3 => n9574, A4 => 
                           n9575, ZN => n9571);
   U13599 : AOI221_X1 port map( B1 => n10650, B2 => n10279, C1 => n10642, C2 =>
                           n9831, A => n9586, ZN => n9569);
   U13600 : AOI221_X1 port map( B1 => n10693, B2 => n10280, C1 => n10685, C2 =>
                           n9832, A => n9585, ZN => n9570);
   U13601 : NOR4_X1 port map( A1 => n9590, A2 => n9591, A3 => n9592, A4 => 
                           n9593, ZN => n9589);
   U13602 : AOI221_X1 port map( B1 => n10650, B2 => n10281, C1 => n10642, C2 =>
                           n9833, A => n9604, ZN => n9587);
   U13603 : AOI221_X1 port map( B1 => n10693, B2 => n10282, C1 => n10685, C2 =>
                           n9834, A => n9603, ZN => n9588);
   U13604 : NOR4_X1 port map( A1 => n9608, A2 => n9609, A3 => n9610, A4 => 
                           n9611, ZN => n9607);
   U13605 : AOI221_X1 port map( B1 => n10650, B2 => n10283, C1 => n10642, C2 =>
                           n9835, A => n9622, ZN => n9605);
   U13606 : AOI221_X1 port map( B1 => n10693, B2 => n10284, C1 => n10685, C2 =>
                           n9836, A => n9621, ZN => n9606);
   U13607 : NOR4_X1 port map( A1 => n9626, A2 => n9627, A3 => n9628, A4 => 
                           n9629, ZN => n9625);
   U13608 : AOI221_X1 port map( B1 => n10650, B2 => n10285, C1 => n10642, C2 =>
                           n9837, A => n9646, ZN => n9623);
   U13609 : AOI221_X1 port map( B1 => n10693, B2 => n10286, C1 => n10685, C2 =>
                           n9838, A => n9644, ZN => n9624);
   U13610 : BUF_X1 port map( A => n7300, Z => n11028);
   U13611 : NOR3_X1 port map( A1 => n6248, A2 => n6249, A3 => n6247, ZN => 
                           n7300);
   U13612 : BUF_X1 port map( A => n8480, Z => n10803);
   U13613 : NOR3_X1 port map( A1 => n6239, A2 => n6240, A3 => n6238, ZN => 
                           n8480);
   U13614 : BUF_X1 port map( A => n11011, Z => n11010);
   U13615 : BUF_X1 port map( A => n11064, Z => n11063);
   U13616 : BUF_X1 port map( A => n11046, Z => n11045);
   U13617 : BUF_X1 port map( A => n10786, Z => n10785);
   U13618 : BUF_X1 port map( A => n10839, Z => n10838);
   U13619 : BUF_X1 port map( A => n10821, Z => n10820);
   U13620 : BUF_X1 port map( A => N2234, Z => n12170);
   U13621 : OAI21_X1 port map( B1 => n7283, B2 => n7286, A => n11507, ZN => 
                           N2234);
   U13622 : BUF_X1 port map( A => N2299, Z => n12161);
   U13623 : OAI21_X1 port map( B1 => n7282, B2 => n7286, A => n11506, ZN => 
                           N2299);
   U13624 : BUF_X1 port map( A => N2364, Z => n12152);
   U13625 : OAI21_X1 port map( B1 => n7281, B2 => n7286, A => n11507, ZN => 
                           N2364);
   U13626 : BUF_X1 port map( A => N2429, Z => n12143);
   U13627 : OAI21_X1 port map( B1 => n7280, B2 => n7286, A => n11506, ZN => 
                           N2429);
   U13628 : BUF_X1 port map( A => N2494, Z => n12134);
   U13629 : OAI21_X1 port map( B1 => n7279, B2 => n7286, A => n11507, ZN => 
                           N2494);
   U13630 : BUF_X1 port map( A => N2559, Z => n12125);
   U13631 : OAI21_X1 port map( B1 => n7278, B2 => n7286, A => n11506, ZN => 
                           N2559);
   U13632 : BUF_X1 port map( A => N2624, Z => n12116);
   U13633 : OAI21_X1 port map( B1 => n7277, B2 => n7286, A => n11508, ZN => 
                           N2624);
   U13634 : BUF_X1 port map( A => N2689, Z => n12107);
   U13635 : OAI21_X1 port map( B1 => n7276, B2 => n7286, A => n11506, ZN => 
                           N2689);
   U13636 : BUF_X1 port map( A => N2754, Z => n12098);
   U13637 : OAI21_X1 port map( B1 => n7283, B2 => n7285, A => n11508, ZN => 
                           N2754);
   U13638 : BUF_X1 port map( A => N2819, Z => n12089);
   U13639 : OAI21_X1 port map( B1 => n7282, B2 => n7285, A => n11506, ZN => 
                           N2819);
   U13640 : BUF_X1 port map( A => N2884, Z => n12080);
   U13641 : OAI21_X1 port map( B1 => n7281, B2 => n7285, A => n11508, ZN => 
                           N2884);
   U13642 : BUF_X1 port map( A => N2949, Z => n12071);
   U13643 : OAI21_X1 port map( B1 => n7280, B2 => n7285, A => n11506, ZN => 
                           N2949);
   U13644 : BUF_X1 port map( A => N3014, Z => n12062);
   U13645 : OAI21_X1 port map( B1 => n7279, B2 => n7285, A => n11507, ZN => 
                           N3014);
   U13646 : BUF_X1 port map( A => N3079, Z => n12053);
   U13647 : OAI21_X1 port map( B1 => n7278, B2 => n7285, A => n11506, ZN => 
                           N3079);
   U13648 : BUF_X1 port map( A => N3144, Z => n12044);
   U13649 : OAI21_X1 port map( B1 => n7277, B2 => n7285, A => n11507, ZN => 
                           N3144);
   U13650 : BUF_X1 port map( A => N3209, Z => n12035);
   U13651 : OAI21_X1 port map( B1 => n7276, B2 => n7285, A => n11507, ZN => 
                           N3209);
   U13652 : BUF_X1 port map( A => N3274, Z => n12026);
   U13653 : OAI21_X1 port map( B1 => n7283, B2 => n7284, A => n11507, ZN => 
                           N3274);
   U13654 : BUF_X1 port map( A => N3339, Z => n12017);
   U13655 : OAI21_X1 port map( B1 => n7282, B2 => n7284, A => n11506, ZN => 
                           N3339);
   U13656 : BUF_X1 port map( A => N3404, Z => n12008);
   U13657 : OAI21_X1 port map( B1 => n7281, B2 => n7284, A => n11508, ZN => 
                           N3404);
   U13658 : BUF_X1 port map( A => N3469, Z => n11999);
   U13659 : OAI21_X1 port map( B1 => n7280, B2 => n7284, A => n11506, ZN => 
                           N3469);
   U13660 : BUF_X1 port map( A => N3534, Z => n11990);
   U13661 : OAI21_X1 port map( B1 => n7279, B2 => n7284, A => n11508, ZN => 
                           N3534);
   U13662 : BUF_X1 port map( A => N3599, Z => n11981);
   U13663 : OAI21_X1 port map( B1 => n7278, B2 => n7284, A => n11506, ZN => 
                           N3599);
   U13664 : BUF_X1 port map( A => N3664, Z => n11972);
   U13665 : OAI21_X1 port map( B1 => n7277, B2 => n7284, A => n11507, ZN => 
                           N3664);
   U13666 : BUF_X1 port map( A => N3729, Z => n11963);
   U13667 : OAI21_X1 port map( B1 => n7276, B2 => n7284, A => n11507, ZN => 
                           N3729);
   U13668 : BUF_X1 port map( A => N3794, Z => n11954);
   U13669 : OAI21_X1 port map( B1 => n7275, B2 => n7283, A => n11507, ZN => 
                           N3794);
   U13670 : BUF_X1 port map( A => N3859, Z => n11945);
   U13671 : OAI21_X1 port map( B1 => n7275, B2 => n7282, A => n11506, ZN => 
                           N3859);
   U13672 : BUF_X1 port map( A => N3924, Z => n11936);
   U13673 : OAI21_X1 port map( B1 => n7275, B2 => n7281, A => n11507, ZN => 
                           N3924);
   U13674 : BUF_X1 port map( A => N3989, Z => n11927);
   U13675 : OAI21_X1 port map( B1 => n7275, B2 => n7280, A => n11506, ZN => 
                           N3989);
   U13676 : BUF_X1 port map( A => N4054, Z => n11918);
   U13677 : OAI21_X1 port map( B1 => n7275, B2 => n7279, A => n11507, ZN => 
                           N4054);
   U13678 : BUF_X1 port map( A => N4119, Z => n11909);
   U13679 : OAI21_X1 port map( B1 => n7275, B2 => n7278, A => n11506, ZN => 
                           N4119);
   U13680 : BUF_X1 port map( A => N4184, Z => n11900);
   U13681 : OAI21_X1 port map( B1 => n7275, B2 => n7277, A => n11507, ZN => 
                           N4184);
   U13682 : BUF_X1 port map( A => n6226, Z => n11882);
   U13683 : BUF_X1 port map( A => n7321, Z => n10883);
   U13684 : NAND2_X1 port map( A1 => n11057, A2 => n8465, ZN => n7321);
   U13685 : BUF_X1 port map( A => n7320, Z => n10892);
   U13686 : NAND2_X1 port map( A1 => n11039, A2 => n8465, ZN => n7320);
   U13687 : BUF_X1 port map( A => n7319, Z => n10901);
   U13688 : NAND2_X1 port map( A1 => n8461, A2 => n8465, ZN => n7319);
   U13689 : BUF_X1 port map( A => n7325, Z => n10858);
   U13690 : NAND2_X1 port map( A1 => n8457, A2 => n8465, ZN => n7325);
   U13691 : BUF_X1 port map( A => n7326, Z => n10849);
   U13692 : NAND2_X1 port map( A1 => n11004, A2 => n8465, ZN => n7326);
   U13693 : BUF_X1 port map( A => n7310, Z => n10959);
   U13694 : NAND2_X1 port map( A1 => n8462, A2 => n8458, ZN => n7310);
   U13695 : BUF_X1 port map( A => n7309, Z => n10968);
   U13696 : NAND2_X1 port map( A1 => n8462, A2 => n8457, ZN => n7309);
   U13697 : BUF_X1 port map( A => n7296, Z => n11065);
   U13698 : NAND2_X1 port map( A1 => n6241, A2 => n6242, ZN => n7296);
   U13699 : BUF_X1 port map( A => n8501, Z => n10658);
   U13700 : NAND2_X1 port map( A1 => n10832, A2 => n9645, ZN => n8501);
   U13701 : BUF_X1 port map( A => n8500, Z => n10667);
   U13702 : NAND2_X1 port map( A1 => n10814, A2 => n9645, ZN => n8500);
   U13703 : BUF_X1 port map( A => n8499, Z => n10676);
   U13704 : NAND2_X1 port map( A1 => n9641, A2 => n9645, ZN => n8499);
   U13705 : BUF_X1 port map( A => n8505, Z => n10633);
   U13706 : NAND2_X1 port map( A1 => n9637, A2 => n9645, ZN => n8505);
   U13707 : BUF_X1 port map( A => n8506, Z => n10624);
   U13708 : NAND2_X1 port map( A1 => n10779, A2 => n9645, ZN => n8506);
   U13709 : BUF_X1 port map( A => n8490, Z => n10734);
   U13710 : NAND2_X1 port map( A1 => n9642, A2 => n9638, ZN => n8490);
   U13711 : BUF_X1 port map( A => n8489, Z => n10743);
   U13712 : NAND2_X1 port map( A1 => n9642, A2 => n9637, ZN => n8489);
   U13713 : BUF_X1 port map( A => n8476, Z => n10840);
   U13714 : NAND2_X1 port map( A1 => n6232, A2 => n6233, ZN => n8476);
   U13715 : INV_X1 port map( A => n8458, ZN => n6246);
   U13716 : INV_X1 port map( A => n8457, ZN => n6245);
   U13717 : INV_X1 port map( A => n8461, ZN => n6243);
   U13718 : INV_X1 port map( A => n8460, ZN => n6244);
   U13719 : INV_X1 port map( A => n9638, ZN => n6237);
   U13720 : INV_X1 port map( A => n9637, ZN => n6236);
   U13721 : INV_X1 port map( A => n9641, ZN => n6234);
   U13722 : INV_X1 port map( A => n9640, ZN => n6235);
   U13723 : BUF_X1 port map( A => n10621, Z => n11530);
   U13724 : BUF_X1 port map( A => n11074, Z => n11075);
   U13725 : BUF_X1 port map( A => n11078, Z => n11079);
   U13726 : BUF_X1 port map( A => n11082, Z => n11083);
   U13727 : BUF_X1 port map( A => n11086, Z => n11087);
   U13728 : BUF_X1 port map( A => n11090, Z => n11091);
   U13729 : BUF_X1 port map( A => n11094, Z => n11095);
   U13730 : BUF_X1 port map( A => n11098, Z => n11099);
   U13731 : BUF_X1 port map( A => n11102, Z => n11103);
   U13732 : BUF_X1 port map( A => n11106, Z => n11107);
   U13733 : BUF_X1 port map( A => n11110, Z => n11111);
   U13734 : BUF_X1 port map( A => n11114, Z => n11115);
   U13735 : BUF_X1 port map( A => n11118, Z => n11119);
   U13736 : BUF_X1 port map( A => n11122, Z => n11123);
   U13737 : BUF_X1 port map( A => n11126, Z => n11127);
   U13738 : BUF_X1 port map( A => n11130, Z => n11131);
   U13739 : BUF_X1 port map( A => n11134, Z => n11135);
   U13740 : BUF_X1 port map( A => n11138, Z => n11139);
   U13741 : BUF_X1 port map( A => n11142, Z => n11143);
   U13742 : BUF_X1 port map( A => n11146, Z => n11147);
   U13743 : BUF_X1 port map( A => n11150, Z => n11151);
   U13744 : BUF_X1 port map( A => n11154, Z => n11155);
   U13745 : BUF_X1 port map( A => n11158, Z => n11159);
   U13746 : BUF_X1 port map( A => n11162, Z => n11163);
   U13747 : BUF_X1 port map( A => n11166, Z => n11167);
   U13748 : BUF_X1 port map( A => n11170, Z => n11171);
   U13749 : BUF_X1 port map( A => n11174, Z => n11175);
   U13750 : BUF_X1 port map( A => n11178, Z => n11179);
   U13751 : BUF_X1 port map( A => n11182, Z => n11183);
   U13752 : BUF_X1 port map( A => n11186, Z => n11187);
   U13753 : BUF_X1 port map( A => n11190, Z => n11191);
   U13754 : BUF_X1 port map( A => n11194, Z => n11195);
   U13755 : BUF_X1 port map( A => n11198, Z => n11199);
   U13756 : BUF_X1 port map( A => n11202, Z => n11203);
   U13757 : BUF_X1 port map( A => n11206, Z => n11207);
   U13758 : BUF_X1 port map( A => n11210, Z => n11211);
   U13759 : BUF_X1 port map( A => n11214, Z => n11215);
   U13760 : BUF_X1 port map( A => n11218, Z => n11219);
   U13761 : BUF_X1 port map( A => n11222, Z => n11223);
   U13762 : BUF_X1 port map( A => n11226, Z => n11227);
   U13763 : BUF_X1 port map( A => n11230, Z => n11231);
   U13764 : BUF_X1 port map( A => n11234, Z => n11235);
   U13765 : BUF_X1 port map( A => n11238, Z => n11239);
   U13766 : BUF_X1 port map( A => n11242, Z => n11243);
   U13767 : BUF_X1 port map( A => n11246, Z => n11247);
   U13768 : BUF_X1 port map( A => n11250, Z => n11251);
   U13769 : BUF_X1 port map( A => n11254, Z => n11255);
   U13770 : BUF_X1 port map( A => n11258, Z => n11259);
   U13771 : BUF_X1 port map( A => n11262, Z => n11263);
   U13772 : BUF_X1 port map( A => n11266, Z => n11267);
   U13773 : BUF_X1 port map( A => n11270, Z => n11271);
   U13774 : BUF_X1 port map( A => n11274, Z => n11275);
   U13775 : BUF_X1 port map( A => n11278, Z => n11279);
   U13776 : BUF_X1 port map( A => n11282, Z => n11283);
   U13777 : BUF_X1 port map( A => n11286, Z => n11287);
   U13778 : BUF_X1 port map( A => n11290, Z => n11291);
   U13779 : BUF_X1 port map( A => n11294, Z => n11295);
   U13780 : BUF_X1 port map( A => n11298, Z => n11299);
   U13781 : BUF_X1 port map( A => n11302, Z => n11303);
   U13782 : BUF_X1 port map( A => n11306, Z => n11307);
   U13783 : BUF_X1 port map( A => n11310, Z => n11311);
   U13784 : BUF_X1 port map( A => n11314, Z => n11315);
   U13785 : BUF_X1 port map( A => n11318, Z => n11319);
   U13786 : BUF_X1 port map( A => n11322, Z => n11323);
   U13787 : BUF_X1 port map( A => n11326, Z => n11327);
   U13788 : BUF_X1 port map( A => n11074, Z => n11076);
   U13789 : BUF_X1 port map( A => n11078, Z => n11080);
   U13790 : BUF_X1 port map( A => n11082, Z => n11084);
   U13791 : BUF_X1 port map( A => n11086, Z => n11088);
   U13792 : BUF_X1 port map( A => n11090, Z => n11092);
   U13793 : BUF_X1 port map( A => n11094, Z => n11096);
   U13794 : BUF_X1 port map( A => n11098, Z => n11100);
   U13795 : BUF_X1 port map( A => n11102, Z => n11104);
   U13796 : BUF_X1 port map( A => n11106, Z => n11108);
   U13797 : BUF_X1 port map( A => n11110, Z => n11112);
   U13798 : BUF_X1 port map( A => n11114, Z => n11116);
   U13799 : BUF_X1 port map( A => n11118, Z => n11120);
   U13800 : BUF_X1 port map( A => n11122, Z => n11124);
   U13801 : BUF_X1 port map( A => n11126, Z => n11128);
   U13802 : BUF_X1 port map( A => n11130, Z => n11132);
   U13803 : BUF_X1 port map( A => n11134, Z => n11136);
   U13804 : BUF_X1 port map( A => n11138, Z => n11140);
   U13805 : BUF_X1 port map( A => n11142, Z => n11144);
   U13806 : BUF_X1 port map( A => n11146, Z => n11148);
   U13807 : BUF_X1 port map( A => n11150, Z => n11152);
   U13808 : BUF_X1 port map( A => n11154, Z => n11156);
   U13809 : BUF_X1 port map( A => n11158, Z => n11160);
   U13810 : BUF_X1 port map( A => n11162, Z => n11164);
   U13811 : BUF_X1 port map( A => n11166, Z => n11168);
   U13812 : BUF_X1 port map( A => n11170, Z => n11172);
   U13813 : BUF_X1 port map( A => n11174, Z => n11176);
   U13814 : BUF_X1 port map( A => n11178, Z => n11180);
   U13815 : BUF_X1 port map( A => n11182, Z => n11184);
   U13816 : BUF_X1 port map( A => n11186, Z => n11188);
   U13817 : BUF_X1 port map( A => n11190, Z => n11192);
   U13818 : BUF_X1 port map( A => n11194, Z => n11196);
   U13819 : BUF_X1 port map( A => n11198, Z => n11200);
   U13820 : BUF_X1 port map( A => n11202, Z => n11204);
   U13821 : BUF_X1 port map( A => n11206, Z => n11208);
   U13822 : BUF_X1 port map( A => n11210, Z => n11212);
   U13823 : BUF_X1 port map( A => n11214, Z => n11216);
   U13824 : BUF_X1 port map( A => n11218, Z => n11220);
   U13825 : BUF_X1 port map( A => n11222, Z => n11224);
   U13826 : BUF_X1 port map( A => n11226, Z => n11228);
   U13827 : BUF_X1 port map( A => n11230, Z => n11232);
   U13828 : BUF_X1 port map( A => n11234, Z => n11236);
   U13829 : BUF_X1 port map( A => n11238, Z => n11240);
   U13830 : BUF_X1 port map( A => n11242, Z => n11244);
   U13831 : BUF_X1 port map( A => n11246, Z => n11248);
   U13832 : BUF_X1 port map( A => n11250, Z => n11252);
   U13833 : BUF_X1 port map( A => n11254, Z => n11256);
   U13834 : BUF_X1 port map( A => n11258, Z => n11260);
   U13835 : BUF_X1 port map( A => n11262, Z => n11264);
   U13836 : BUF_X1 port map( A => n11266, Z => n11268);
   U13837 : BUF_X1 port map( A => n11270, Z => n11272);
   U13838 : BUF_X1 port map( A => n11274, Z => n11276);
   U13839 : BUF_X1 port map( A => n11278, Z => n11280);
   U13840 : BUF_X1 port map( A => n11282, Z => n11284);
   U13841 : BUF_X1 port map( A => n11286, Z => n11288);
   U13842 : BUF_X1 port map( A => n11290, Z => n11292);
   U13843 : BUF_X1 port map( A => n11294, Z => n11296);
   U13844 : BUF_X1 port map( A => n11298, Z => n11300);
   U13845 : BUF_X1 port map( A => n11302, Z => n11304);
   U13846 : BUF_X1 port map( A => n11306, Z => n11308);
   U13847 : BUF_X1 port map( A => n11310, Z => n11312);
   U13848 : BUF_X1 port map( A => n11314, Z => n11316);
   U13849 : BUF_X1 port map( A => n11318, Z => n11320);
   U13850 : BUF_X1 port map( A => n11322, Z => n11324);
   U13851 : BUF_X1 port map( A => n11326, Z => n11328);
   U13852 : BUF_X1 port map( A => n11074, Z => n11077);
   U13853 : BUF_X1 port map( A => n11078, Z => n11081);
   U13854 : BUF_X1 port map( A => n11082, Z => n11085);
   U13855 : BUF_X1 port map( A => n11086, Z => n11089);
   U13856 : BUF_X1 port map( A => n11090, Z => n11093);
   U13857 : BUF_X1 port map( A => n11094, Z => n11097);
   U13858 : BUF_X1 port map( A => n11098, Z => n11101);
   U13859 : BUF_X1 port map( A => n11102, Z => n11105);
   U13860 : BUF_X1 port map( A => n11106, Z => n11109);
   U13861 : BUF_X1 port map( A => n11110, Z => n11113);
   U13862 : BUF_X1 port map( A => n11114, Z => n11117);
   U13863 : BUF_X1 port map( A => n11118, Z => n11121);
   U13864 : BUF_X1 port map( A => n11122, Z => n11125);
   U13865 : BUF_X1 port map( A => n11126, Z => n11129);
   U13866 : BUF_X1 port map( A => n11130, Z => n11133);
   U13867 : BUF_X1 port map( A => n11134, Z => n11137);
   U13868 : BUF_X1 port map( A => n11138, Z => n11141);
   U13869 : BUF_X1 port map( A => n11142, Z => n11145);
   U13870 : BUF_X1 port map( A => n11146, Z => n11149);
   U13871 : BUF_X1 port map( A => n11150, Z => n11153);
   U13872 : BUF_X1 port map( A => n11154, Z => n11157);
   U13873 : BUF_X1 port map( A => n11158, Z => n11161);
   U13874 : BUF_X1 port map( A => n11162, Z => n11165);
   U13875 : BUF_X1 port map( A => n11166, Z => n11169);
   U13876 : BUF_X1 port map( A => n11170, Z => n11173);
   U13877 : BUF_X1 port map( A => n11174, Z => n11177);
   U13878 : BUF_X1 port map( A => n11178, Z => n11181);
   U13879 : BUF_X1 port map( A => n11182, Z => n11185);
   U13880 : BUF_X1 port map( A => n11186, Z => n11189);
   U13881 : BUF_X1 port map( A => n11190, Z => n11193);
   U13882 : BUF_X1 port map( A => n11194, Z => n11197);
   U13883 : BUF_X1 port map( A => n11198, Z => n11201);
   U13884 : BUF_X1 port map( A => n11202, Z => n11205);
   U13885 : BUF_X1 port map( A => n11206, Z => n11209);
   U13886 : BUF_X1 port map( A => n11210, Z => n11213);
   U13887 : BUF_X1 port map( A => n11214, Z => n11217);
   U13888 : BUF_X1 port map( A => n11218, Z => n11221);
   U13889 : BUF_X1 port map( A => n11222, Z => n11225);
   U13890 : BUF_X1 port map( A => n11226, Z => n11229);
   U13891 : BUF_X1 port map( A => n11230, Z => n11233);
   U13892 : BUF_X1 port map( A => n11234, Z => n11237);
   U13893 : BUF_X1 port map( A => n11238, Z => n11241);
   U13894 : BUF_X1 port map( A => n11242, Z => n11245);
   U13895 : BUF_X1 port map( A => n11246, Z => n11249);
   U13896 : BUF_X1 port map( A => n11250, Z => n11253);
   U13897 : BUF_X1 port map( A => n11254, Z => n11257);
   U13898 : BUF_X1 port map( A => n11258, Z => n11261);
   U13899 : BUF_X1 port map( A => n11262, Z => n11265);
   U13900 : BUF_X1 port map( A => n11266, Z => n11269);
   U13901 : BUF_X1 port map( A => n11270, Z => n11273);
   U13902 : BUF_X1 port map( A => n11274, Z => n11277);
   U13903 : BUF_X1 port map( A => n11278, Z => n11281);
   U13904 : BUF_X1 port map( A => n11282, Z => n11285);
   U13905 : BUF_X1 port map( A => n11286, Z => n11289);
   U13906 : BUF_X1 port map( A => n11290, Z => n11293);
   U13907 : BUF_X1 port map( A => n11294, Z => n11297);
   U13908 : BUF_X1 port map( A => n11298, Z => n11301);
   U13909 : BUF_X1 port map( A => n11302, Z => n11305);
   U13910 : BUF_X1 port map( A => n11306, Z => n11309);
   U13911 : BUF_X1 port map( A => n11310, Z => n11313);
   U13912 : BUF_X1 port map( A => n11314, Z => n11317);
   U13913 : BUF_X1 port map( A => n11318, Z => n11321);
   U13914 : BUF_X1 port map( A => n11322, Z => n11325);
   U13915 : BUF_X1 port map( A => n11326, Z => n11329);
   U13916 : NOR2_X1 port map( A1 => n6241, A2 => ADD_RD2(3), ZN => n8465);
   U13917 : NOR2_X1 port map( A1 => n6232, A2 => ADD_RD1(3), ZN => n9645);
   U13918 : NOR3_X1 port map( A1 => n6248, A2 => ADD_RD2(0), A3 => n6247, ZN =>
                           n8457);
   U13919 : NOR3_X1 port map( A1 => n6239, A2 => ADD_RD1(0), A3 => n6238, ZN =>
                           n9637);
   U13920 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n6247, 
                           ZN => n8458);
   U13921 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n6238, 
                           ZN => n9638);
   U13922 : OAI222_X1 port map( A1 => n1152_port, A2 => n10907, B1 => 
                           n1088_port, B2 => n10898, C1 => n1216_port, C2 => 
                           n10889, ZN => n7318);
   U13923 : OAI222_X1 port map( A1 => n1151_port, A2 => n10907, B1 => 
                           n1087_port, B2 => n10898, C1 => n1215_port, C2 => 
                           n10889, ZN => n7343);
   U13924 : OAI222_X1 port map( A1 => n1150_port, A2 => n10907, B1 => 
                           n1086_port, B2 => n10898, C1 => n1214_port, C2 => 
                           n10889, ZN => n7361);
   U13925 : OAI222_X1 port map( A1 => n1149_port, A2 => n10907, B1 => 
                           n1085_port, B2 => n10898, C1 => n1213_port, C2 => 
                           n10889, ZN => n7379);
   U13926 : OAI222_X1 port map( A1 => n1148_port, A2 => n10906, B1 => 
                           n1084_port, B2 => n10897, C1 => n1212_port, C2 => 
                           n10888, ZN => n7397);
   U13927 : OAI222_X1 port map( A1 => n1147_port, A2 => n10906, B1 => 
                           n1083_port, B2 => n10897, C1 => n1211_port, C2 => 
                           n10888, ZN => n7415);
   U13928 : OAI222_X1 port map( A1 => n1146_port, A2 => n10906, B1 => 
                           n1082_port, B2 => n10897, C1 => n1210_port, C2 => 
                           n10888, ZN => n7433);
   U13929 : OAI222_X1 port map( A1 => n1145_port, A2 => n10906, B1 => 
                           n1081_port, B2 => n10897, C1 => n1209_port, C2 => 
                           n10888, ZN => n7451);
   U13930 : OAI222_X1 port map( A1 => n1144_port, A2 => n10906, B1 => 
                           n1080_port, B2 => n10897, C1 => n1208_port, C2 => 
                           n10888, ZN => n7469);
   U13931 : OAI222_X1 port map( A1 => n1143_port, A2 => n10906, B1 => 
                           n1079_port, B2 => n10897, C1 => n1207_port, C2 => 
                           n10888, ZN => n7487);
   U13932 : OAI222_X1 port map( A1 => n1142_port, A2 => n10906, B1 => 
                           n1078_port, B2 => n10897, C1 => n1206_port, C2 => 
                           n10888, ZN => n7505);
   U13933 : OAI222_X1 port map( A1 => n1141_port, A2 => n10906, B1 => 
                           n1077_port, B2 => n10897, C1 => n1205_port, C2 => 
                           n10888, ZN => n7523);
   U13934 : OAI222_X1 port map( A1 => n1140_port, A2 => n10906, B1 => 
                           n1076_port, B2 => n10897, C1 => n1204_port, C2 => 
                           n10888, ZN => n7541);
   U13935 : OAI222_X1 port map( A1 => n1139_port, A2 => n10906, B1 => 
                           n1075_port, B2 => n10897, C1 => n1203_port, C2 => 
                           n10888, ZN => n7559);
   U13936 : OAI222_X1 port map( A1 => n1138_port, A2 => n10906, B1 => 
                           n1074_port, B2 => n10897, C1 => n1202_port, C2 => 
                           n10888, ZN => n7577);
   U13937 : OAI222_X1 port map( A1 => n1137_port, A2 => n10906, B1 => 
                           n1073_port, B2 => n10897, C1 => n1201_port, C2 => 
                           n10888, ZN => n7595);
   U13938 : OAI222_X1 port map( A1 => n1136_port, A2 => n10905, B1 => 
                           n1072_port, B2 => n10896, C1 => n1200_port, C2 => 
                           n10887, ZN => n7613);
   U13939 : OAI222_X1 port map( A1 => n1135_port, A2 => n10905, B1 => 
                           n1071_port, B2 => n10896, C1 => n1199_port, C2 => 
                           n10887, ZN => n7631);
   U13940 : OAI222_X1 port map( A1 => n1134_port, A2 => n10905, B1 => 
                           n1070_port, B2 => n10896, C1 => n1198_port, C2 => 
                           n10887, ZN => n7649);
   U13941 : OAI222_X1 port map( A1 => n1133_port, A2 => n10905, B1 => 
                           n1069_port, B2 => n10896, C1 => n1197_port, C2 => 
                           n10887, ZN => n7667);
   U13942 : OAI222_X1 port map( A1 => n1132_port, A2 => n10905, B1 => 
                           n1068_port, B2 => n10896, C1 => n1196_port, C2 => 
                           n10887, ZN => n7685);
   U13943 : OAI222_X1 port map( A1 => n1131_port, A2 => n10905, B1 => 
                           n1067_port, B2 => n10896, C1 => n1195_port, C2 => 
                           n10887, ZN => n7703);
   U13944 : OAI222_X1 port map( A1 => n1130_port, A2 => n10905, B1 => 
                           n1066_port, B2 => n10896, C1 => n1194_port, C2 => 
                           n10887, ZN => n7721);
   U13945 : OAI222_X1 port map( A1 => n1129_port, A2 => n10905, B1 => 
                           n1065_port, B2 => n10896, C1 => n1193_port, C2 => 
                           n10887, ZN => n7739);
   U13946 : OAI222_X1 port map( A1 => n1128_port, A2 => n10905, B1 => 
                           n1064_port, B2 => n10896, C1 => n1192_port, C2 => 
                           n10887, ZN => n7757);
   U13947 : OAI222_X1 port map( A1 => n1127_port, A2 => n10905, B1 => 
                           n1063_port, B2 => n10896, C1 => n1191_port, C2 => 
                           n10887, ZN => n7775);
   U13948 : OAI222_X1 port map( A1 => n1126_port, A2 => n10905, B1 => 
                           n1062_port, B2 => n10896, C1 => n1190_port, C2 => 
                           n10887, ZN => n7793);
   U13949 : OAI222_X1 port map( A1 => n1125_port, A2 => n10905, B1 => 
                           n1061_port, B2 => n10896, C1 => n1189_port, C2 => 
                           n10887, ZN => n7811);
   U13950 : OAI222_X1 port map( A1 => n1124_port, A2 => n10904, B1 => 
                           n1060_port, B2 => n10895, C1 => n1188_port, C2 => 
                           n10886, ZN => n7829);
   U13951 : OAI222_X1 port map( A1 => n1123_port, A2 => n10904, B1 => 
                           n1059_port, B2 => n10895, C1 => n1187_port, C2 => 
                           n10886, ZN => n7847);
   U13952 : OAI222_X1 port map( A1 => n1122_port, A2 => n10904, B1 => 
                           n1058_port, B2 => n10895, C1 => n1186_port, C2 => 
                           n10886, ZN => n7865);
   U13953 : OAI222_X1 port map( A1 => n1121_port, A2 => n10904, B1 => 
                           n1057_port, B2 => n10895, C1 => n1185_port, C2 => 
                           n10886, ZN => n7883);
   U13954 : OAI222_X1 port map( A1 => n1120_port, A2 => n10904, B1 => 
                           n1056_port, B2 => n10895, C1 => n1184_port, C2 => 
                           n10886, ZN => n7901);
   U13955 : OAI222_X1 port map( A1 => n1119_port, A2 => n10904, B1 => 
                           n1055_port, B2 => n10895, C1 => n1183_port, C2 => 
                           n10886, ZN => n7919);
   U13956 : OAI222_X1 port map( A1 => n1118_port, A2 => n10904, B1 => 
                           n1054_port, B2 => n10895, C1 => n1182_port, C2 => 
                           n10886, ZN => n7937);
   U13957 : OAI222_X1 port map( A1 => n1117_port, A2 => n10904, B1 => 
                           n1053_port, B2 => n10895, C1 => n1181_port, C2 => 
                           n10886, ZN => n7955);
   U13958 : OAI222_X1 port map( A1 => n1116_port, A2 => n10904, B1 => 
                           n1052_port, B2 => n10895, C1 => n1180_port, C2 => 
                           n10886, ZN => n7973);
   U13959 : OAI222_X1 port map( A1 => n1115_port, A2 => n10904, B1 => 
                           n1051_port, B2 => n10895, C1 => n1179_port, C2 => 
                           n10886, ZN => n7991);
   U13960 : OAI222_X1 port map( A1 => n1114_port, A2 => n10904, B1 => 
                           n1050_port, B2 => n10895, C1 => n1178_port, C2 => 
                           n10886, ZN => n8009);
   U13961 : OAI222_X1 port map( A1 => n1113_port, A2 => n10904, B1 => 
                           n1049_port, B2 => n10895, C1 => n1177_port, C2 => 
                           n10886, ZN => n8027);
   U13962 : OAI222_X1 port map( A1 => n1112_port, A2 => n10903, B1 => 
                           n1048_port, B2 => n10894, C1 => n1176_port, C2 => 
                           n10885, ZN => n8045);
   U13963 : OAI222_X1 port map( A1 => n1111_port, A2 => n10903, B1 => 
                           n1047_port, B2 => n10894, C1 => n1175_port, C2 => 
                           n10885, ZN => n8063);
   U13964 : OAI222_X1 port map( A1 => n1110_port, A2 => n10903, B1 => 
                           n1046_port, B2 => n10894, C1 => n1174_port, C2 => 
                           n10885, ZN => n8081);
   U13965 : OAI222_X1 port map( A1 => n1109_port, A2 => n10903, B1 => 
                           n1045_port, B2 => n10894, C1 => n1173_port, C2 => 
                           n10885, ZN => n8099);
   U13966 : OAI222_X1 port map( A1 => n1108_port, A2 => n10903, B1 => 
                           n1044_port, B2 => n10894, C1 => n1172_port, C2 => 
                           n10885, ZN => n8117);
   U13967 : OAI222_X1 port map( A1 => n1107_port, A2 => n10903, B1 => 
                           n1043_port, B2 => n10894, C1 => n1171_port, C2 => 
                           n10885, ZN => n8135);
   U13968 : OAI222_X1 port map( A1 => n1106_port, A2 => n10903, B1 => 
                           n1042_port, B2 => n10894, C1 => n1170_port, C2 => 
                           n10885, ZN => n8153);
   U13969 : OAI222_X1 port map( A1 => n1105_port, A2 => n10903, B1 => 
                           n1041_port, B2 => n10894, C1 => n1169_port, C2 => 
                           n10885, ZN => n8171);
   U13970 : OAI222_X1 port map( A1 => n1104_port, A2 => n10903, B1 => 
                           n1040_port, B2 => n10894, C1 => n1168_port, C2 => 
                           n10885, ZN => n8189);
   U13971 : OAI222_X1 port map( A1 => n1103_port, A2 => n10903, B1 => 
                           n1039_port, B2 => n10894, C1 => n1167_port, C2 => 
                           n10885, ZN => n8207);
   U13972 : OAI222_X1 port map( A1 => n1102_port, A2 => n10903, B1 => 
                           n1038_port, B2 => n10894, C1 => n1166_port, C2 => 
                           n10885, ZN => n8225);
   U13973 : OAI222_X1 port map( A1 => n1101_port, A2 => n10903, B1 => 
                           n1037_port, B2 => n10894, C1 => n1165_port, C2 => 
                           n10885, ZN => n8243);
   U13974 : OAI222_X1 port map( A1 => n1100_port, A2 => n10902, B1 => 
                           n1036_port, B2 => n10893, C1 => n1164_port, C2 => 
                           n10884, ZN => n8261);
   U13975 : OAI222_X1 port map( A1 => n1099_port, A2 => n10902, B1 => 
                           n1035_port, B2 => n10893, C1 => n1163_port, C2 => 
                           n10884, ZN => n8279);
   U13976 : OAI222_X1 port map( A1 => n1098_port, A2 => n10902, B1 => 
                           n1034_port, B2 => n10893, C1 => n1162_port, C2 => 
                           n10884, ZN => n8297);
   U13977 : OAI222_X1 port map( A1 => n1097_port, A2 => n10902, B1 => 
                           n1033_port, B2 => n10893, C1 => n1161_port, C2 => 
                           n10884, ZN => n8315);
   U13978 : OAI222_X1 port map( A1 => n1096_port, A2 => n10902, B1 => 
                           n1032_port, B2 => n10893, C1 => n1160_port, C2 => 
                           n10884, ZN => n8333);
   U13979 : OAI222_X1 port map( A1 => n1095_port, A2 => n10902, B1 => 
                           n1031_port, B2 => n10893, C1 => n1159_port, C2 => 
                           n10884, ZN => n8351);
   U13980 : OAI222_X1 port map( A1 => n1094_port, A2 => n10902, B1 => 
                           n1030_port, B2 => n10893, C1 => n1158_port, C2 => 
                           n10884, ZN => n8369);
   U13981 : OAI222_X1 port map( A1 => n1093_port, A2 => n10902, B1 => 
                           n1029_port, B2 => n10893, C1 => n1157_port, C2 => 
                           n10884, ZN => n8387);
   U13982 : OAI222_X1 port map( A1 => n1092_port, A2 => n10902, B1 => 
                           n1028_port, B2 => n10893, C1 => n1156_port, C2 => 
                           n10884, ZN => n8405);
   U13983 : OAI222_X1 port map( A1 => n1091_port, A2 => n10902, B1 => 
                           n1027_port, B2 => n10893, C1 => n1155_port, C2 => 
                           n10884, ZN => n8423);
   U13984 : OAI222_X1 port map( A1 => n1090_port, A2 => n10902, B1 => 
                           n1026_port, B2 => n10893, C1 => n1154_port, C2 => 
                           n10884, ZN => n8441);
   U13985 : OAI222_X1 port map( A1 => n1089_port, A2 => n10902, B1 => 
                           n1025_port, B2 => n10893, C1 => n1153_port, C2 => 
                           n10884, ZN => n8464);
   U13986 : OAI222_X1 port map( A1 => n1152_port, A2 => n10682, B1 => 
                           n1088_port, B2 => n10673, C1 => n1216_port, C2 => 
                           n10664, ZN => n8498);
   U13987 : OAI222_X1 port map( A1 => n1151_port, A2 => n10682, B1 => 
                           n1087_port, B2 => n10673, C1 => n1215_port, C2 => 
                           n10664, ZN => n8523);
   U13988 : OAI222_X1 port map( A1 => n1150_port, A2 => n10682, B1 => 
                           n1086_port, B2 => n10673, C1 => n1214_port, C2 => 
                           n10664, ZN => n8541);
   U13989 : OAI222_X1 port map( A1 => n1149_port, A2 => n10682, B1 => 
                           n1085_port, B2 => n10673, C1 => n1213_port, C2 => 
                           n10664, ZN => n8559);
   U13990 : OAI222_X1 port map( A1 => n1148_port, A2 => n10681, B1 => 
                           n1084_port, B2 => n10672, C1 => n1212_port, C2 => 
                           n10663, ZN => n8577);
   U13991 : OAI222_X1 port map( A1 => n1147_port, A2 => n10681, B1 => 
                           n1083_port, B2 => n10672, C1 => n1211_port, C2 => 
                           n10663, ZN => n8595);
   U13992 : OAI222_X1 port map( A1 => n1146_port, A2 => n10681, B1 => 
                           n1082_port, B2 => n10672, C1 => n1210_port, C2 => 
                           n10663, ZN => n8613);
   U13993 : OAI222_X1 port map( A1 => n1145_port, A2 => n10681, B1 => 
                           n1081_port, B2 => n10672, C1 => n1209_port, C2 => 
                           n10663, ZN => n8631);
   U13994 : OAI222_X1 port map( A1 => n1144_port, A2 => n10681, B1 => 
                           n1080_port, B2 => n10672, C1 => n1208_port, C2 => 
                           n10663, ZN => n8649);
   U13995 : OAI222_X1 port map( A1 => n1143_port, A2 => n10681, B1 => 
                           n1079_port, B2 => n10672, C1 => n1207_port, C2 => 
                           n10663, ZN => n8667);
   U13996 : OAI222_X1 port map( A1 => n1142_port, A2 => n10681, B1 => 
                           n1078_port, B2 => n10672, C1 => n1206_port, C2 => 
                           n10663, ZN => n8685);
   U13997 : OAI222_X1 port map( A1 => n1141_port, A2 => n10681, B1 => 
                           n1077_port, B2 => n10672, C1 => n1205_port, C2 => 
                           n10663, ZN => n8703);
   U13998 : OAI222_X1 port map( A1 => n1140_port, A2 => n10681, B1 => 
                           n1076_port, B2 => n10672, C1 => n1204_port, C2 => 
                           n10663, ZN => n8721);
   U13999 : OAI222_X1 port map( A1 => n1139_port, A2 => n10681, B1 => 
                           n1075_port, B2 => n10672, C1 => n1203_port, C2 => 
                           n10663, ZN => n8739);
   U14000 : OAI222_X1 port map( A1 => n1138_port, A2 => n10681, B1 => 
                           n1074_port, B2 => n10672, C1 => n1202_port, C2 => 
                           n10663, ZN => n8757);
   U14001 : OAI222_X1 port map( A1 => n1137_port, A2 => n10681, B1 => 
                           n1073_port, B2 => n10672, C1 => n1201_port, C2 => 
                           n10663, ZN => n8775);
   U14002 : OAI222_X1 port map( A1 => n1136_port, A2 => n10680, B1 => 
                           n1072_port, B2 => n10671, C1 => n1200_port, C2 => 
                           n10662, ZN => n8793);
   U14003 : OAI222_X1 port map( A1 => n1135_port, A2 => n10680, B1 => 
                           n1071_port, B2 => n10671, C1 => n1199_port, C2 => 
                           n10662, ZN => n8811);
   U14004 : OAI222_X1 port map( A1 => n1134_port, A2 => n10680, B1 => 
                           n1070_port, B2 => n10671, C1 => n1198_port, C2 => 
                           n10662, ZN => n8829);
   U14005 : OAI222_X1 port map( A1 => n1133_port, A2 => n10680, B1 => 
                           n1069_port, B2 => n10671, C1 => n1197_port, C2 => 
                           n10662, ZN => n8847);
   U14006 : OAI222_X1 port map( A1 => n1132_port, A2 => n10680, B1 => 
                           n1068_port, B2 => n10671, C1 => n1196_port, C2 => 
                           n10662, ZN => n8865);
   U14007 : OAI222_X1 port map( A1 => n1131_port, A2 => n10680, B1 => 
                           n1067_port, B2 => n10671, C1 => n1195_port, C2 => 
                           n10662, ZN => n8883);
   U14008 : OAI222_X1 port map( A1 => n1130_port, A2 => n10680, B1 => 
                           n1066_port, B2 => n10671, C1 => n1194_port, C2 => 
                           n10662, ZN => n8901);
   U14009 : OAI222_X1 port map( A1 => n1129_port, A2 => n10680, B1 => 
                           n1065_port, B2 => n10671, C1 => n1193_port, C2 => 
                           n10662, ZN => n8919);
   U14010 : OAI222_X1 port map( A1 => n1128_port, A2 => n10680, B1 => 
                           n1064_port, B2 => n10671, C1 => n1192_port, C2 => 
                           n10662, ZN => n8937);
   U14011 : OAI222_X1 port map( A1 => n1127_port, A2 => n10680, B1 => 
                           n1063_port, B2 => n10671, C1 => n1191_port, C2 => 
                           n10662, ZN => n8955);
   U14012 : OAI222_X1 port map( A1 => n1126_port, A2 => n10680, B1 => 
                           n1062_port, B2 => n10671, C1 => n1190_port, C2 => 
                           n10662, ZN => n8973);
   U14013 : OAI222_X1 port map( A1 => n1125_port, A2 => n10680, B1 => 
                           n1061_port, B2 => n10671, C1 => n1189_port, C2 => 
                           n10662, ZN => n8991);
   U14014 : OAI222_X1 port map( A1 => n1124_port, A2 => n10679, B1 => 
                           n1060_port, B2 => n10670, C1 => n1188_port, C2 => 
                           n10661, ZN => n9009);
   U14015 : OAI222_X1 port map( A1 => n1123_port, A2 => n10679, B1 => 
                           n1059_port, B2 => n10670, C1 => n1187_port, C2 => 
                           n10661, ZN => n9027);
   U14016 : OAI222_X1 port map( A1 => n1122_port, A2 => n10679, B1 => 
                           n1058_port, B2 => n10670, C1 => n1186_port, C2 => 
                           n10661, ZN => n9045);
   U14017 : OAI222_X1 port map( A1 => n1121_port, A2 => n10679, B1 => 
                           n1057_port, B2 => n10670, C1 => n1185_port, C2 => 
                           n10661, ZN => n9063);
   U14018 : OAI222_X1 port map( A1 => n1120_port, A2 => n10679, B1 => 
                           n1056_port, B2 => n10670, C1 => n1184_port, C2 => 
                           n10661, ZN => n9081);
   U14019 : OAI222_X1 port map( A1 => n1119_port, A2 => n10679, B1 => 
                           n1055_port, B2 => n10670, C1 => n1183_port, C2 => 
                           n10661, ZN => n9099);
   U14020 : OAI222_X1 port map( A1 => n1118_port, A2 => n10679, B1 => 
                           n1054_port, B2 => n10670, C1 => n1182_port, C2 => 
                           n10661, ZN => n9117);
   U14021 : OAI222_X1 port map( A1 => n1117_port, A2 => n10679, B1 => 
                           n1053_port, B2 => n10670, C1 => n1181_port, C2 => 
                           n10661, ZN => n9135);
   U14022 : OAI222_X1 port map( A1 => n1116_port, A2 => n10679, B1 => 
                           n1052_port, B2 => n10670, C1 => n1180_port, C2 => 
                           n10661, ZN => n9153);
   U14023 : OAI222_X1 port map( A1 => n1115_port, A2 => n10679, B1 => 
                           n1051_port, B2 => n10670, C1 => n1179_port, C2 => 
                           n10661, ZN => n9171);
   U14024 : OAI222_X1 port map( A1 => n1114_port, A2 => n10679, B1 => 
                           n1050_port, B2 => n10670, C1 => n1178_port, C2 => 
                           n10661, ZN => n9189);
   U14025 : OAI222_X1 port map( A1 => n1113_port, A2 => n10679, B1 => 
                           n1049_port, B2 => n10670, C1 => n1177_port, C2 => 
                           n10661, ZN => n9207);
   U14026 : OAI222_X1 port map( A1 => n1112_port, A2 => n10678, B1 => 
                           n1048_port, B2 => n10669, C1 => n1176_port, C2 => 
                           n10660, ZN => n9225);
   U14027 : OAI222_X1 port map( A1 => n1111_port, A2 => n10678, B1 => 
                           n1047_port, B2 => n10669, C1 => n1175_port, C2 => 
                           n10660, ZN => n9243);
   U14028 : OAI222_X1 port map( A1 => n1110_port, A2 => n10678, B1 => 
                           n1046_port, B2 => n10669, C1 => n1174_port, C2 => 
                           n10660, ZN => n9261);
   U14029 : OAI222_X1 port map( A1 => n1109_port, A2 => n10678, B1 => 
                           n1045_port, B2 => n10669, C1 => n1173_port, C2 => 
                           n10660, ZN => n9279);
   U14030 : OAI222_X1 port map( A1 => n1108_port, A2 => n10678, B1 => 
                           n1044_port, B2 => n10669, C1 => n1172_port, C2 => 
                           n10660, ZN => n9297);
   U14031 : OAI222_X1 port map( A1 => n1107_port, A2 => n10678, B1 => 
                           n1043_port, B2 => n10669, C1 => n1171_port, C2 => 
                           n10660, ZN => n9315);
   U14032 : OAI222_X1 port map( A1 => n1106_port, A2 => n10678, B1 => 
                           n1042_port, B2 => n10669, C1 => n1170_port, C2 => 
                           n10660, ZN => n9333);
   U14033 : OAI222_X1 port map( A1 => n1105_port, A2 => n10678, B1 => 
                           n1041_port, B2 => n10669, C1 => n1169_port, C2 => 
                           n10660, ZN => n9351);
   U14034 : OAI222_X1 port map( A1 => n1104_port, A2 => n10678, B1 => 
                           n1040_port, B2 => n10669, C1 => n1168_port, C2 => 
                           n10660, ZN => n9369);
   U14035 : OAI222_X1 port map( A1 => n1103_port, A2 => n10678, B1 => 
                           n1039_port, B2 => n10669, C1 => n1167_port, C2 => 
                           n10660, ZN => n9387);
   U14036 : OAI222_X1 port map( A1 => n1102_port, A2 => n10678, B1 => 
                           n1038_port, B2 => n10669, C1 => n1166_port, C2 => 
                           n10660, ZN => n9405);
   U14037 : OAI222_X1 port map( A1 => n1101_port, A2 => n10678, B1 => 
                           n1037_port, B2 => n10669, C1 => n1165_port, C2 => 
                           n10660, ZN => n9423);
   U14038 : OAI222_X1 port map( A1 => n1100_port, A2 => n10677, B1 => 
                           n1036_port, B2 => n10668, C1 => n1164_port, C2 => 
                           n10659, ZN => n9441);
   U14039 : OAI222_X1 port map( A1 => n1099_port, A2 => n10677, B1 => 
                           n1035_port, B2 => n10668, C1 => n1163_port, C2 => 
                           n10659, ZN => n9459);
   U14040 : OAI222_X1 port map( A1 => n1098_port, A2 => n10677, B1 => 
                           n1034_port, B2 => n10668, C1 => n1162_port, C2 => 
                           n10659, ZN => n9477);
   U14041 : OAI222_X1 port map( A1 => n1097_port, A2 => n10677, B1 => 
                           n1033_port, B2 => n10668, C1 => n1161_port, C2 => 
                           n10659, ZN => n9495);
   U14042 : OAI222_X1 port map( A1 => n1096_port, A2 => n10677, B1 => 
                           n1032_port, B2 => n10668, C1 => n1160_port, C2 => 
                           n10659, ZN => n9513);
   U14043 : OAI222_X1 port map( A1 => n1095_port, A2 => n10677, B1 => 
                           n1031_port, B2 => n10668, C1 => n1159_port, C2 => 
                           n10659, ZN => n9531);
   U14044 : OAI222_X1 port map( A1 => n1094_port, A2 => n10677, B1 => 
                           n1030_port, B2 => n10668, C1 => n1158_port, C2 => 
                           n10659, ZN => n9549);
   U14045 : OAI222_X1 port map( A1 => n1093_port, A2 => n10677, B1 => 
                           n1029_port, B2 => n10668, C1 => n1157_port, C2 => 
                           n10659, ZN => n9567);
   U14046 : OAI222_X1 port map( A1 => n1092_port, A2 => n10677, B1 => 
                           n1028_port, B2 => n10668, C1 => n1156_port, C2 => 
                           n10659, ZN => n9585);
   U14047 : OAI222_X1 port map( A1 => n1091_port, A2 => n10677, B1 => 
                           n1027_port, B2 => n10668, C1 => n1155_port, C2 => 
                           n10659, ZN => n9603);
   U14048 : OAI222_X1 port map( A1 => n1090_port, A2 => n10677, B1 => 
                           n1026_port, B2 => n10668, C1 => n1154_port, C2 => 
                           n10659, ZN => n9621);
   U14049 : OAI222_X1 port map( A1 => n1089_port, A2 => n10677, B1 => 
                           n1025_port, B2 => n10668, C1 => n1153_port, C2 => 
                           n10659, ZN => n9644);
   U14050 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n6249, 
                           ZN => n8461);
   U14051 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n6240, 
                           ZN => n9641);
   U14052 : NOR3_X1 port map( A1 => n6249, A2 => ADD_RD2(2), A3 => n6248, ZN =>
                           n8460);
   U14053 : NOR3_X1 port map( A1 => n6240, A2 => ADD_RD1(2), A3 => n6239, ZN =>
                           n9640);
   U14054 : NAND2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n7286);
   U14055 : NAND2_X1 port map( A1 => ADD_WR(4), A2 => n6228, ZN => n7285);
   U14056 : NAND2_X1 port map( A1 => ADD_WR(3), A2 => n6227, ZN => n7284);
   U14057 : OAI221_X1 port map( B1 => n1856_port, B2 => n10965, C1 => 
                           n1920_port, C2 => n10956, A => n7312, ZN => n7290);
   U14058 : AOI222_X1 port map( A1 => n10947, A2 => n9647, B1 => n10939, B2 => 
                           n10095, C1 => n10931, C2 => n10543, ZN => n7312);
   U14059 : OAI221_X1 port map( B1 => n1855_port, B2 => n10965, C1 => 
                           n1919_port, C2 => n10956, A => n7342, ZN => n7330);
   U14060 : AOI222_X1 port map( A1 => n10947, A2 => n9648, B1 => n10939, B2 => 
                           n10096, C1 => n10931, C2 => n10544, ZN => n7342);
   U14061 : OAI221_X1 port map( B1 => n1854_port, B2 => n10965, C1 => 
                           n1918_port, C2 => n10956, A => n7360, ZN => n7348);
   U14062 : AOI222_X1 port map( A1 => n10947, A2 => n9649, B1 => n10939, B2 => 
                           n10097, C1 => n10931, C2 => n10545, ZN => n7360);
   U14063 : OAI221_X1 port map( B1 => n1853_port, B2 => n10965, C1 => 
                           n1917_port, C2 => n10956, A => n7378, ZN => n7366);
   U14064 : AOI222_X1 port map( A1 => n10947, A2 => n9650, B1 => n10939, B2 => 
                           n10098, C1 => n10931, C2 => n10546, ZN => n7378);
   U14065 : OAI221_X1 port map( B1 => n1852_port, B2 => n10964, C1 => 
                           n1916_port, C2 => n10955, A => n7396, ZN => n7384);
   U14066 : AOI222_X1 port map( A1 => n10946, A2 => n9651, B1 => n10938, B2 => 
                           n10099, C1 => n10930, C2 => n10547, ZN => n7396);
   U14067 : OAI221_X1 port map( B1 => n1851_port, B2 => n10964, C1 => 
                           n1915_port, C2 => n10955, A => n7414, ZN => n7402);
   U14068 : AOI222_X1 port map( A1 => n10946, A2 => n9652, B1 => n10938, B2 => 
                           n10100, C1 => n10930, C2 => n10548, ZN => n7414);
   U14069 : OAI221_X1 port map( B1 => n1850_port, B2 => n10964, C1 => 
                           n1914_port, C2 => n10955, A => n7432, ZN => n7420);
   U14070 : AOI222_X1 port map( A1 => n10946, A2 => n9653, B1 => n10938, B2 => 
                           n10101, C1 => n10930, C2 => n10549, ZN => n7432);
   U14071 : OAI221_X1 port map( B1 => n1849_port, B2 => n10964, C1 => 
                           n1913_port, C2 => n10955, A => n7450, ZN => n7438);
   U14072 : AOI222_X1 port map( A1 => n10946, A2 => n9654, B1 => n10938, B2 => 
                           n10102, C1 => n10930, C2 => n10550, ZN => n7450);
   U14073 : OAI221_X1 port map( B1 => n1848_port, B2 => n10964, C1 => 
                           n1912_port, C2 => n10955, A => n7468, ZN => n7456);
   U14074 : AOI222_X1 port map( A1 => n10946, A2 => n9655, B1 => n10938, B2 => 
                           n10103, C1 => n10930, C2 => n10551, ZN => n7468);
   U14075 : OAI221_X1 port map( B1 => n1847_port, B2 => n10964, C1 => 
                           n1911_port, C2 => n10955, A => n7486, ZN => n7474);
   U14076 : AOI222_X1 port map( A1 => n10946, A2 => n9656, B1 => n10938, B2 => 
                           n10104, C1 => n10930, C2 => n10552, ZN => n7486);
   U14077 : OAI221_X1 port map( B1 => n1846_port, B2 => n10964, C1 => 
                           n1910_port, C2 => n10955, A => n7504, ZN => n7492);
   U14078 : AOI222_X1 port map( A1 => n10946, A2 => n9657, B1 => n10938, B2 => 
                           n10105, C1 => n10930, C2 => n10553, ZN => n7504);
   U14079 : OAI221_X1 port map( B1 => n1845_port, B2 => n10964, C1 => 
                           n1909_port, C2 => n10955, A => n7522, ZN => n7510);
   U14080 : AOI222_X1 port map( A1 => n10946, A2 => n9658, B1 => n10938, B2 => 
                           n10106, C1 => n10930, C2 => n10554, ZN => n7522);
   U14081 : OAI221_X1 port map( B1 => n1844_port, B2 => n10964, C1 => 
                           n1908_port, C2 => n10955, A => n7540, ZN => n7528);
   U14082 : AOI222_X1 port map( A1 => n10946, A2 => n9659, B1 => n10938, B2 => 
                           n10107, C1 => n10930, C2 => n10555, ZN => n7540);
   U14083 : OAI221_X1 port map( B1 => n1843_port, B2 => n10964, C1 => 
                           n1907_port, C2 => n10955, A => n7558, ZN => n7546);
   U14084 : AOI222_X1 port map( A1 => n10946, A2 => n9660, B1 => n10938, B2 => 
                           n10108, C1 => n10930, C2 => n10556, ZN => n7558);
   U14085 : OAI221_X1 port map( B1 => n1842_port, B2 => n10964, C1 => 
                           n1906_port, C2 => n10955, A => n7576, ZN => n7564);
   U14086 : AOI222_X1 port map( A1 => n10946, A2 => n9661, B1 => n10938, B2 => 
                           n10109, C1 => n10930, C2 => n10557, ZN => n7576);
   U14087 : OAI221_X1 port map( B1 => n1841_port, B2 => n10964, C1 => 
                           n1905_port, C2 => n10955, A => n7594, ZN => n7582);
   U14088 : AOI222_X1 port map( A1 => n10946, A2 => n9662, B1 => n10938, B2 => 
                           n10110, C1 => n10930, C2 => n10558, ZN => n7594);
   U14089 : OAI221_X1 port map( B1 => n1840_port, B2 => n10963, C1 => 
                           n1904_port, C2 => n10954, A => n7612, ZN => n7600);
   U14090 : AOI222_X1 port map( A1 => n10945, A2 => n9663, B1 => n10937, B2 => 
                           n10111, C1 => n10929, C2 => n10559, ZN => n7612);
   U14091 : OAI221_X1 port map( B1 => n1839_port, B2 => n10963, C1 => 
                           n1903_port, C2 => n10954, A => n7630, ZN => n7618);
   U14092 : AOI222_X1 port map( A1 => n10945, A2 => n9664, B1 => n10937, B2 => 
                           n10112, C1 => n10929, C2 => n10560, ZN => n7630);
   U14093 : OAI221_X1 port map( B1 => n1838_port, B2 => n10963, C1 => 
                           n1902_port, C2 => n10954, A => n7648, ZN => n7636);
   U14094 : AOI222_X1 port map( A1 => n10945, A2 => n9665, B1 => n10937, B2 => 
                           n10113, C1 => n10929, C2 => n10561, ZN => n7648);
   U14095 : OAI221_X1 port map( B1 => n1837_port, B2 => n10963, C1 => 
                           n1901_port, C2 => n10954, A => n7666, ZN => n7654);
   U14096 : AOI222_X1 port map( A1 => n10945, A2 => n9666, B1 => n10937, B2 => 
                           n10114, C1 => n10929, C2 => n10562, ZN => n7666);
   U14097 : OAI221_X1 port map( B1 => n1836_port, B2 => n10963, C1 => 
                           n1900_port, C2 => n10954, A => n7684, ZN => n7672);
   U14098 : AOI222_X1 port map( A1 => n10945, A2 => n9667, B1 => n10937, B2 => 
                           n10115, C1 => n10929, C2 => n10563, ZN => n7684);
   U14099 : OAI221_X1 port map( B1 => n1835_port, B2 => n10963, C1 => 
                           n1899_port, C2 => n10954, A => n7702, ZN => n7690);
   U14100 : AOI222_X1 port map( A1 => n10945, A2 => n9668, B1 => n10937, B2 => 
                           n10116, C1 => n10929, C2 => n10564, ZN => n7702);
   U14101 : OAI221_X1 port map( B1 => n1834_port, B2 => n10963, C1 => 
                           n1898_port, C2 => n10954, A => n7720, ZN => n7708);
   U14102 : AOI222_X1 port map( A1 => n10945, A2 => n9669, B1 => n10937, B2 => 
                           n10117, C1 => n10929, C2 => n10565, ZN => n7720);
   U14103 : OAI221_X1 port map( B1 => n1833_port, B2 => n10963, C1 => 
                           n1897_port, C2 => n10954, A => n7738, ZN => n7726);
   U14104 : AOI222_X1 port map( A1 => n10945, A2 => n9670, B1 => n10937, B2 => 
                           n10118, C1 => n10929, C2 => n10566, ZN => n7738);
   U14105 : OAI221_X1 port map( B1 => n1832_port, B2 => n10963, C1 => 
                           n1896_port, C2 => n10954, A => n7756, ZN => n7744);
   U14106 : AOI222_X1 port map( A1 => n10945, A2 => n9671, B1 => n10937, B2 => 
                           n10119, C1 => n10929, C2 => n10567, ZN => n7756);
   U14107 : OAI221_X1 port map( B1 => n1831_port, B2 => n10963, C1 => 
                           n1895_port, C2 => n10954, A => n7774, ZN => n7762);
   U14108 : AOI222_X1 port map( A1 => n10945, A2 => n9672, B1 => n10937, B2 => 
                           n10120, C1 => n10929, C2 => n10568, ZN => n7774);
   U14109 : OAI221_X1 port map( B1 => n1830_port, B2 => n10963, C1 => 
                           n1894_port, C2 => n10954, A => n7792, ZN => n7780);
   U14110 : AOI222_X1 port map( A1 => n10945, A2 => n9673, B1 => n10937, B2 => 
                           n10121, C1 => n10929, C2 => n10569, ZN => n7792);
   U14111 : OAI221_X1 port map( B1 => n1829_port, B2 => n10963, C1 => 
                           n1893_port, C2 => n10954, A => n7810, ZN => n7798);
   U14112 : AOI222_X1 port map( A1 => n10945, A2 => n9674, B1 => n10937, B2 => 
                           n10122, C1 => n10929, C2 => n10570, ZN => n7810);
   U14113 : OAI221_X1 port map( B1 => n1828_port, B2 => n10962, C1 => 
                           n1892_port, C2 => n10953, A => n7828, ZN => n7816);
   U14114 : AOI222_X1 port map( A1 => n10944, A2 => n9675, B1 => n10936, B2 => 
                           n10123, C1 => n10928, C2 => n10571, ZN => n7828);
   U14115 : OAI221_X1 port map( B1 => n1827_port, B2 => n10962, C1 => 
                           n1891_port, C2 => n10953, A => n7846, ZN => n7834);
   U14116 : AOI222_X1 port map( A1 => n10944, A2 => n9676, B1 => n10936, B2 => 
                           n10124, C1 => n10928, C2 => n10572, ZN => n7846);
   U14117 : OAI221_X1 port map( B1 => n1826_port, B2 => n10962, C1 => 
                           n1890_port, C2 => n10953, A => n7864, ZN => n7852);
   U14118 : AOI222_X1 port map( A1 => n10944, A2 => n9677, B1 => n10936, B2 => 
                           n10125, C1 => n10928, C2 => n10573, ZN => n7864);
   U14119 : OAI221_X1 port map( B1 => n1825_port, B2 => n10962, C1 => 
                           n1889_port, C2 => n10953, A => n7882, ZN => n7870);
   U14120 : AOI222_X1 port map( A1 => n10944, A2 => n9678, B1 => n10936, B2 => 
                           n10126, C1 => n10928, C2 => n10574, ZN => n7882);
   U14121 : OAI221_X1 port map( B1 => n1824_port, B2 => n10962, C1 => 
                           n1888_port, C2 => n10953, A => n7900, ZN => n7888);
   U14122 : AOI222_X1 port map( A1 => n10944, A2 => n9679, B1 => n10936, B2 => 
                           n10127, C1 => n10928, C2 => n10575, ZN => n7900);
   U14123 : OAI221_X1 port map( B1 => n1823_port, B2 => n10962, C1 => 
                           n1887_port, C2 => n10953, A => n7918, ZN => n7906);
   U14124 : AOI222_X1 port map( A1 => n10944, A2 => n9680, B1 => n10936, B2 => 
                           n10128, C1 => n10928, C2 => n10576, ZN => n7918);
   U14125 : OAI221_X1 port map( B1 => n1822_port, B2 => n10962, C1 => 
                           n1886_port, C2 => n10953, A => n7936, ZN => n7924);
   U14126 : AOI222_X1 port map( A1 => n10944, A2 => n9681, B1 => n10936, B2 => 
                           n10129, C1 => n10928, C2 => n10577, ZN => n7936);
   U14127 : OAI221_X1 port map( B1 => n1821_port, B2 => n10962, C1 => 
                           n1885_port, C2 => n10953, A => n7954, ZN => n7942);
   U14128 : AOI222_X1 port map( A1 => n10944, A2 => n9682, B1 => n10936, B2 => 
                           n10130, C1 => n10928, C2 => n10578, ZN => n7954);
   U14129 : OAI221_X1 port map( B1 => n1820_port, B2 => n10962, C1 => 
                           n1884_port, C2 => n10953, A => n7972, ZN => n7960);
   U14130 : AOI222_X1 port map( A1 => n10944, A2 => n9683, B1 => n10936, B2 => 
                           n10131, C1 => n10928, C2 => n10579, ZN => n7972);
   U14131 : OAI221_X1 port map( B1 => n1819_port, B2 => n10962, C1 => 
                           n1883_port, C2 => n10953, A => n7990, ZN => n7978);
   U14132 : AOI222_X1 port map( A1 => n10944, A2 => n9684, B1 => n10936, B2 => 
                           n10132, C1 => n10928, C2 => n10580, ZN => n7990);
   U14133 : OAI221_X1 port map( B1 => n1818_port, B2 => n10962, C1 => 
                           n1882_port, C2 => n10953, A => n8008, ZN => n7996);
   U14134 : AOI222_X1 port map( A1 => n10944, A2 => n9685, B1 => n10936, B2 => 
                           n10133, C1 => n10928, C2 => n10581, ZN => n8008);
   U14135 : OAI221_X1 port map( B1 => n1817_port, B2 => n10962, C1 => 
                           n1881_port, C2 => n10953, A => n8026, ZN => n8014);
   U14136 : AOI222_X1 port map( A1 => n10944, A2 => n9686, B1 => n10936, B2 => 
                           n10134, C1 => n10928, C2 => n10582, ZN => n8026);
   U14137 : OAI221_X1 port map( B1 => n1816_port, B2 => n10961, C1 => 
                           n1880_port, C2 => n10952, A => n8044, ZN => n8032);
   U14138 : AOI222_X1 port map( A1 => n10943, A2 => n9687, B1 => n10935, B2 => 
                           n10135, C1 => n10927, C2 => n10583, ZN => n8044);
   U14139 : OAI221_X1 port map( B1 => n1815_port, B2 => n10961, C1 => 
                           n1879_port, C2 => n10952, A => n8062, ZN => n8050);
   U14140 : AOI222_X1 port map( A1 => n10943, A2 => n9688, B1 => n10935, B2 => 
                           n10136, C1 => n10927, C2 => n10584, ZN => n8062);
   U14141 : OAI221_X1 port map( B1 => n1814_port, B2 => n10961, C1 => 
                           n1878_port, C2 => n10952, A => n8080, ZN => n8068);
   U14142 : AOI222_X1 port map( A1 => n10943, A2 => n9689, B1 => n10935, B2 => 
                           n10137, C1 => n10927, C2 => n10585, ZN => n8080);
   U14143 : OAI221_X1 port map( B1 => n1813_port, B2 => n10961, C1 => 
                           n1877_port, C2 => n10952, A => n8098, ZN => n8086);
   U14144 : AOI222_X1 port map( A1 => n10943, A2 => n9690, B1 => n10935, B2 => 
                           n10138, C1 => n10927, C2 => n10586, ZN => n8098);
   U14145 : OAI221_X1 port map( B1 => n1812_port, B2 => n10961, C1 => 
                           n1876_port, C2 => n10952, A => n8116, ZN => n8104);
   U14146 : AOI222_X1 port map( A1 => n10943, A2 => n9691, B1 => n10935, B2 => 
                           n10139, C1 => n10927, C2 => n10587, ZN => n8116);
   U14147 : OAI221_X1 port map( B1 => n1811_port, B2 => n10961, C1 => 
                           n1875_port, C2 => n10952, A => n8134, ZN => n8122);
   U14148 : AOI222_X1 port map( A1 => n10943, A2 => n9692, B1 => n10935, B2 => 
                           n10140, C1 => n10927, C2 => n10588, ZN => n8134);
   U14149 : OAI221_X1 port map( B1 => n1810_port, B2 => n10961, C1 => 
                           n1874_port, C2 => n10952, A => n8152, ZN => n8140);
   U14150 : AOI222_X1 port map( A1 => n10943, A2 => n9693, B1 => n10935, B2 => 
                           n10141, C1 => n10927, C2 => n10589, ZN => n8152);
   U14151 : OAI221_X1 port map( B1 => n1809_port, B2 => n10961, C1 => 
                           n1873_port, C2 => n10952, A => n8170, ZN => n8158);
   U14152 : AOI222_X1 port map( A1 => n10943, A2 => n9694, B1 => n10935, B2 => 
                           n10142, C1 => n10927, C2 => n10590, ZN => n8170);
   U14153 : OAI221_X1 port map( B1 => n1808_port, B2 => n10961, C1 => 
                           n1872_port, C2 => n10952, A => n8188, ZN => n8176);
   U14154 : AOI222_X1 port map( A1 => n10943, A2 => n9695, B1 => n10935, B2 => 
                           n10143, C1 => n10927, C2 => n10591, ZN => n8188);
   U14155 : OAI221_X1 port map( B1 => n1807_port, B2 => n10961, C1 => 
                           n1871_port, C2 => n10952, A => n8206, ZN => n8194);
   U14156 : AOI222_X1 port map( A1 => n10943, A2 => n9696, B1 => n10935, B2 => 
                           n10144, C1 => n10927, C2 => n10592, ZN => n8206);
   U14157 : OAI221_X1 port map( B1 => n1806_port, B2 => n10961, C1 => 
                           n1870_port, C2 => n10952, A => n8224, ZN => n8212);
   U14158 : AOI222_X1 port map( A1 => n10943, A2 => n9697, B1 => n10935, B2 => 
                           n10145, C1 => n10927, C2 => n10593, ZN => n8224);
   U14159 : OAI221_X1 port map( B1 => n1805_port, B2 => n10961, C1 => 
                           n1869_port, C2 => n10952, A => n8242, ZN => n8230);
   U14160 : AOI222_X1 port map( A1 => n10943, A2 => n9698, B1 => n10935, B2 => 
                           n10146, C1 => n10927, C2 => n10594, ZN => n8242);
   U14161 : OAI221_X1 port map( B1 => n1804_port, B2 => n10960, C1 => 
                           n1868_port, C2 => n10951, A => n8260, ZN => n8248);
   U14162 : AOI222_X1 port map( A1 => n10942, A2 => n9699, B1 => n10934, B2 => 
                           n10147, C1 => n10926, C2 => n10595, ZN => n8260);
   U14163 : OAI221_X1 port map( B1 => n1803_port, B2 => n10960, C1 => 
                           n1867_port, C2 => n10951, A => n8278, ZN => n8266);
   U14164 : AOI222_X1 port map( A1 => n10942, A2 => n9700, B1 => n10934, B2 => 
                           n10148, C1 => n10926, C2 => n10596, ZN => n8278);
   U14165 : OAI221_X1 port map( B1 => n1802_port, B2 => n10960, C1 => 
                           n1866_port, C2 => n10951, A => n8296, ZN => n8284);
   U14166 : AOI222_X1 port map( A1 => n10942, A2 => n9701, B1 => n10934, B2 => 
                           n10149, C1 => n10926, C2 => n10597, ZN => n8296);
   U14167 : OAI221_X1 port map( B1 => n1801_port, B2 => n10960, C1 => 
                           n1865_port, C2 => n10951, A => n8314, ZN => n8302);
   U14168 : AOI222_X1 port map( A1 => n10942, A2 => n9702, B1 => n10934, B2 => 
                           n10150, C1 => n10926, C2 => n10598, ZN => n8314);
   U14169 : OAI221_X1 port map( B1 => n1800_port, B2 => n10960, C1 => 
                           n1864_port, C2 => n10951, A => n8332, ZN => n8320);
   U14170 : AOI222_X1 port map( A1 => n10942, A2 => n9703, B1 => n10934, B2 => 
                           n10151, C1 => n10926, C2 => n10599, ZN => n8332);
   U14171 : OAI221_X1 port map( B1 => n1799_port, B2 => n10960, C1 => 
                           n1863_port, C2 => n10951, A => n8350, ZN => n8338);
   U14172 : AOI222_X1 port map( A1 => n10942, A2 => n9704, B1 => n10934, B2 => 
                           n10152, C1 => n10926, C2 => n10600, ZN => n8350);
   U14173 : OAI221_X1 port map( B1 => n1798_port, B2 => n10960, C1 => 
                           n1862_port, C2 => n10951, A => n8368, ZN => n8356);
   U14174 : AOI222_X1 port map( A1 => n10942, A2 => n9705, B1 => n10934, B2 => 
                           n10153, C1 => n10926, C2 => n10601, ZN => n8368);
   U14175 : OAI221_X1 port map( B1 => n1797_port, B2 => n10960, C1 => 
                           n1861_port, C2 => n10951, A => n8386, ZN => n8374);
   U14176 : AOI222_X1 port map( A1 => n10942, A2 => n9706, B1 => n10934, B2 => 
                           n10154, C1 => n10926, C2 => n10602, ZN => n8386);
   U14177 : OAI221_X1 port map( B1 => n1796_port, B2 => n10960, C1 => 
                           n1860_port, C2 => n10951, A => n8404, ZN => n8392);
   U14178 : AOI222_X1 port map( A1 => n10942, A2 => n9707, B1 => n10934, B2 => 
                           n10155, C1 => n10926, C2 => n10603, ZN => n8404);
   U14179 : OAI221_X1 port map( B1 => n1795_port, B2 => n10960, C1 => 
                           n1859_port, C2 => n10951, A => n8422, ZN => n8410);
   U14180 : AOI222_X1 port map( A1 => n10942, A2 => n9708, B1 => n10934, B2 => 
                           n10156, C1 => n10926, C2 => n10604, ZN => n8422);
   U14181 : OAI221_X1 port map( B1 => n1794_port, B2 => n10960, C1 => 
                           n1858_port, C2 => n10951, A => n8440, ZN => n8428);
   U14182 : AOI222_X1 port map( A1 => n10942, A2 => n9709, B1 => n10934, B2 => 
                           n10157, C1 => n10926, C2 => n10605, ZN => n8440);
   U14183 : OAI221_X1 port map( B1 => n1793_port, B2 => n10960, C1 => 
                           n1857_port, C2 => n10951, A => n8463, ZN => n8446);
   U14184 : AOI222_X1 port map( A1 => n10942, A2 => n9710, B1 => n10934, B2 => 
                           n10158, C1 => n10926, C2 => n10606, ZN => n8463);
   U14185 : OAI221_X1 port map( B1 => n1856_port, B2 => n10740, C1 => 
                           n1920_port, C2 => n10731, A => n8492, ZN => n8470);
   U14186 : AOI222_X1 port map( A1 => n10722, A2 => n9647, B1 => n10714, B2 => 
                           n10095, C1 => n10706, C2 => n10543, ZN => n8492);
   U14187 : OAI221_X1 port map( B1 => n1855_port, B2 => n10740, C1 => 
                           n1919_port, C2 => n10731, A => n8522, ZN => n8510);
   U14188 : AOI222_X1 port map( A1 => n10722, A2 => n9648, B1 => n10714, B2 => 
                           n10096, C1 => n10706, C2 => n10544, ZN => n8522);
   U14189 : OAI221_X1 port map( B1 => n1854_port, B2 => n10740, C1 => 
                           n1918_port, C2 => n10731, A => n8540, ZN => n8528);
   U14190 : AOI222_X1 port map( A1 => n10722, A2 => n9649, B1 => n10714, B2 => 
                           n10097, C1 => n10706, C2 => n10545, ZN => n8540);
   U14191 : OAI221_X1 port map( B1 => n1853_port, B2 => n10740, C1 => 
                           n1917_port, C2 => n10731, A => n8558, ZN => n8546);
   U14192 : AOI222_X1 port map( A1 => n10722, A2 => n9650, B1 => n10714, B2 => 
                           n10098, C1 => n10706, C2 => n10546, ZN => n8558);
   U14193 : OAI221_X1 port map( B1 => n1852_port, B2 => n10739, C1 => 
                           n1916_port, C2 => n10730, A => n8576, ZN => n8564);
   U14194 : AOI222_X1 port map( A1 => n10721, A2 => n9651, B1 => n10713, B2 => 
                           n10099, C1 => n10705, C2 => n10547, ZN => n8576);
   U14195 : OAI221_X1 port map( B1 => n1851_port, B2 => n10739, C1 => 
                           n1915_port, C2 => n10730, A => n8594, ZN => n8582);
   U14196 : AOI222_X1 port map( A1 => n10721, A2 => n9652, B1 => n10713, B2 => 
                           n10100, C1 => n10705, C2 => n10548, ZN => n8594);
   U14197 : OAI221_X1 port map( B1 => n1850_port, B2 => n10739, C1 => 
                           n1914_port, C2 => n10730, A => n8612, ZN => n8600);
   U14198 : AOI222_X1 port map( A1 => n10721, A2 => n9653, B1 => n10713, B2 => 
                           n10101, C1 => n10705, C2 => n10549, ZN => n8612);
   U14199 : OAI221_X1 port map( B1 => n1849_port, B2 => n10739, C1 => 
                           n1913_port, C2 => n10730, A => n8630, ZN => n8618);
   U14200 : AOI222_X1 port map( A1 => n10721, A2 => n9654, B1 => n10713, B2 => 
                           n10102, C1 => n10705, C2 => n10550, ZN => n8630);
   U14201 : OAI221_X1 port map( B1 => n1848_port, B2 => n10739, C1 => 
                           n1912_port, C2 => n10730, A => n8648, ZN => n8636);
   U14202 : AOI222_X1 port map( A1 => n10721, A2 => n9655, B1 => n10713, B2 => 
                           n10103, C1 => n10705, C2 => n10551, ZN => n8648);
   U14203 : OAI221_X1 port map( B1 => n1847_port, B2 => n10739, C1 => 
                           n1911_port, C2 => n10730, A => n8666, ZN => n8654);
   U14204 : AOI222_X1 port map( A1 => n10721, A2 => n9656, B1 => n10713, B2 => 
                           n10104, C1 => n10705, C2 => n10552, ZN => n8666);
   U14205 : OAI221_X1 port map( B1 => n1846_port, B2 => n10739, C1 => 
                           n1910_port, C2 => n10730, A => n8684, ZN => n8672);
   U14206 : AOI222_X1 port map( A1 => n10721, A2 => n9657, B1 => n10713, B2 => 
                           n10105, C1 => n10705, C2 => n10553, ZN => n8684);
   U14207 : OAI221_X1 port map( B1 => n1845_port, B2 => n10739, C1 => 
                           n1909_port, C2 => n10730, A => n8702, ZN => n8690);
   U14208 : AOI222_X1 port map( A1 => n10721, A2 => n9658, B1 => n10713, B2 => 
                           n10106, C1 => n10705, C2 => n10554, ZN => n8702);
   U14209 : OAI221_X1 port map( B1 => n1844_port, B2 => n10739, C1 => 
                           n1908_port, C2 => n10730, A => n8720, ZN => n8708);
   U14210 : AOI222_X1 port map( A1 => n10721, A2 => n9659, B1 => n10713, B2 => 
                           n10107, C1 => n10705, C2 => n10555, ZN => n8720);
   U14211 : OAI221_X1 port map( B1 => n1843_port, B2 => n10739, C1 => 
                           n1907_port, C2 => n10730, A => n8738, ZN => n8726);
   U14212 : AOI222_X1 port map( A1 => n10721, A2 => n9660, B1 => n10713, B2 => 
                           n10108, C1 => n10705, C2 => n10556, ZN => n8738);
   U14213 : OAI221_X1 port map( B1 => n1842_port, B2 => n10739, C1 => 
                           n1906_port, C2 => n10730, A => n8756, ZN => n8744);
   U14214 : AOI222_X1 port map( A1 => n10721, A2 => n9661, B1 => n10713, B2 => 
                           n10109, C1 => n10705, C2 => n10557, ZN => n8756);
   U14215 : OAI221_X1 port map( B1 => n1841_port, B2 => n10739, C1 => 
                           n1905_port, C2 => n10730, A => n8774, ZN => n8762);
   U14216 : AOI222_X1 port map( A1 => n10721, A2 => n9662, B1 => n10713, B2 => 
                           n10110, C1 => n10705, C2 => n10558, ZN => n8774);
   U14217 : OAI221_X1 port map( B1 => n1840_port, B2 => n10738, C1 => 
                           n1904_port, C2 => n10729, A => n8792, ZN => n8780);
   U14218 : AOI222_X1 port map( A1 => n10720, A2 => n9663, B1 => n10712, B2 => 
                           n10111, C1 => n10704, C2 => n10559, ZN => n8792);
   U14219 : OAI221_X1 port map( B1 => n1839_port, B2 => n10738, C1 => 
                           n1903_port, C2 => n10729, A => n8810, ZN => n8798);
   U14220 : AOI222_X1 port map( A1 => n10720, A2 => n9664, B1 => n10712, B2 => 
                           n10112, C1 => n10704, C2 => n10560, ZN => n8810);
   U14221 : OAI221_X1 port map( B1 => n1838_port, B2 => n10738, C1 => 
                           n1902_port, C2 => n10729, A => n8828, ZN => n8816);
   U14222 : AOI222_X1 port map( A1 => n10720, A2 => n9665, B1 => n10712, B2 => 
                           n10113, C1 => n10704, C2 => n10561, ZN => n8828);
   U14223 : OAI221_X1 port map( B1 => n1837_port, B2 => n10738, C1 => 
                           n1901_port, C2 => n10729, A => n8846, ZN => n8834);
   U14224 : AOI222_X1 port map( A1 => n10720, A2 => n9666, B1 => n10712, B2 => 
                           n10114, C1 => n10704, C2 => n10562, ZN => n8846);
   U14225 : OAI221_X1 port map( B1 => n1836_port, B2 => n10738, C1 => 
                           n1900_port, C2 => n10729, A => n8864, ZN => n8852);
   U14226 : AOI222_X1 port map( A1 => n10720, A2 => n9667, B1 => n10712, B2 => 
                           n10115, C1 => n10704, C2 => n10563, ZN => n8864);
   U14227 : OAI221_X1 port map( B1 => n1835_port, B2 => n10738, C1 => 
                           n1899_port, C2 => n10729, A => n8882, ZN => n8870);
   U14228 : AOI222_X1 port map( A1 => n10720, A2 => n9668, B1 => n10712, B2 => 
                           n10116, C1 => n10704, C2 => n10564, ZN => n8882);
   U14229 : OAI221_X1 port map( B1 => n1834_port, B2 => n10738, C1 => 
                           n1898_port, C2 => n10729, A => n8900, ZN => n8888);
   U14230 : AOI222_X1 port map( A1 => n10720, A2 => n9669, B1 => n10712, B2 => 
                           n10117, C1 => n10704, C2 => n10565, ZN => n8900);
   U14231 : OAI221_X1 port map( B1 => n1833_port, B2 => n10738, C1 => 
                           n1897_port, C2 => n10729, A => n8918, ZN => n8906);
   U14232 : AOI222_X1 port map( A1 => n10720, A2 => n9670, B1 => n10712, B2 => 
                           n10118, C1 => n10704, C2 => n10566, ZN => n8918);
   U14233 : OAI221_X1 port map( B1 => n1832_port, B2 => n10738, C1 => 
                           n1896_port, C2 => n10729, A => n8936, ZN => n8924);
   U14234 : AOI222_X1 port map( A1 => n10720, A2 => n9671, B1 => n10712, B2 => 
                           n10119, C1 => n10704, C2 => n10567, ZN => n8936);
   U14235 : OAI221_X1 port map( B1 => n1831_port, B2 => n10738, C1 => 
                           n1895_port, C2 => n10729, A => n8954, ZN => n8942);
   U14236 : AOI222_X1 port map( A1 => n10720, A2 => n9672, B1 => n10712, B2 => 
                           n10120, C1 => n10704, C2 => n10568, ZN => n8954);
   U14237 : OAI221_X1 port map( B1 => n1830_port, B2 => n10738, C1 => 
                           n1894_port, C2 => n10729, A => n8972, ZN => n8960);
   U14238 : AOI222_X1 port map( A1 => n10720, A2 => n9673, B1 => n10712, B2 => 
                           n10121, C1 => n10704, C2 => n10569, ZN => n8972);
   U14239 : OAI221_X1 port map( B1 => n1829_port, B2 => n10738, C1 => 
                           n1893_port, C2 => n10729, A => n8990, ZN => n8978);
   U14240 : AOI222_X1 port map( A1 => n10720, A2 => n9674, B1 => n10712, B2 => 
                           n10122, C1 => n10704, C2 => n10570, ZN => n8990);
   U14241 : OAI221_X1 port map( B1 => n1828_port, B2 => n10737, C1 => 
                           n1892_port, C2 => n10728, A => n9008, ZN => n8996);
   U14242 : AOI222_X1 port map( A1 => n10719, A2 => n9675, B1 => n10711, B2 => 
                           n10123, C1 => n10703, C2 => n10571, ZN => n9008);
   U14243 : OAI221_X1 port map( B1 => n1827_port, B2 => n10737, C1 => 
                           n1891_port, C2 => n10728, A => n9026, ZN => n9014);
   U14244 : AOI222_X1 port map( A1 => n10719, A2 => n9676, B1 => n10711, B2 => 
                           n10124, C1 => n10703, C2 => n10572, ZN => n9026);
   U14245 : OAI221_X1 port map( B1 => n1826_port, B2 => n10737, C1 => 
                           n1890_port, C2 => n10728, A => n9044, ZN => n9032);
   U14246 : AOI222_X1 port map( A1 => n10719, A2 => n9677, B1 => n10711, B2 => 
                           n10125, C1 => n10703, C2 => n10573, ZN => n9044);
   U14247 : OAI221_X1 port map( B1 => n1825_port, B2 => n10737, C1 => 
                           n1889_port, C2 => n10728, A => n9062, ZN => n9050);
   U14248 : AOI222_X1 port map( A1 => n10719, A2 => n9678, B1 => n10711, B2 => 
                           n10126, C1 => n10703, C2 => n10574, ZN => n9062);
   U14249 : OAI221_X1 port map( B1 => n1824_port, B2 => n10737, C1 => 
                           n1888_port, C2 => n10728, A => n9080, ZN => n9068);
   U14250 : AOI222_X1 port map( A1 => n10719, A2 => n9679, B1 => n10711, B2 => 
                           n10127, C1 => n10703, C2 => n10575, ZN => n9080);
   U14251 : OAI221_X1 port map( B1 => n1823_port, B2 => n10737, C1 => 
                           n1887_port, C2 => n10728, A => n9098, ZN => n9086);
   U14252 : AOI222_X1 port map( A1 => n10719, A2 => n9680, B1 => n10711, B2 => 
                           n10128, C1 => n10703, C2 => n10576, ZN => n9098);
   U14253 : OAI221_X1 port map( B1 => n1822_port, B2 => n10737, C1 => 
                           n1886_port, C2 => n10728, A => n9116, ZN => n9104);
   U14254 : AOI222_X1 port map( A1 => n10719, A2 => n9681, B1 => n10711, B2 => 
                           n10129, C1 => n10703, C2 => n10577, ZN => n9116);
   U14255 : OAI221_X1 port map( B1 => n1821_port, B2 => n10737, C1 => 
                           n1885_port, C2 => n10728, A => n9134, ZN => n9122);
   U14256 : AOI222_X1 port map( A1 => n10719, A2 => n9682, B1 => n10711, B2 => 
                           n10130, C1 => n10703, C2 => n10578, ZN => n9134);
   U14257 : OAI221_X1 port map( B1 => n1820_port, B2 => n10737, C1 => 
                           n1884_port, C2 => n10728, A => n9152, ZN => n9140);
   U14258 : AOI222_X1 port map( A1 => n10719, A2 => n9683, B1 => n10711, B2 => 
                           n10131, C1 => n10703, C2 => n10579, ZN => n9152);
   U14259 : OAI221_X1 port map( B1 => n1819_port, B2 => n10737, C1 => 
                           n1883_port, C2 => n10728, A => n9170, ZN => n9158);
   U14260 : AOI222_X1 port map( A1 => n10719, A2 => n9684, B1 => n10711, B2 => 
                           n10132, C1 => n10703, C2 => n10580, ZN => n9170);
   U14261 : OAI221_X1 port map( B1 => n1818_port, B2 => n10737, C1 => 
                           n1882_port, C2 => n10728, A => n9188, ZN => n9176);
   U14262 : AOI222_X1 port map( A1 => n10719, A2 => n9685, B1 => n10711, B2 => 
                           n10133, C1 => n10703, C2 => n10581, ZN => n9188);
   U14263 : OAI221_X1 port map( B1 => n1817_port, B2 => n10737, C1 => 
                           n1881_port, C2 => n10728, A => n9206, ZN => n9194);
   U14264 : AOI222_X1 port map( A1 => n10719, A2 => n9686, B1 => n10711, B2 => 
                           n10134, C1 => n10703, C2 => n10582, ZN => n9206);
   U14265 : OAI221_X1 port map( B1 => n1816_port, B2 => n10736, C1 => 
                           n1880_port, C2 => n10727, A => n9224, ZN => n9212);
   U14266 : AOI222_X1 port map( A1 => n10718, A2 => n9687, B1 => n10710, B2 => 
                           n10135, C1 => n10702, C2 => n10583, ZN => n9224);
   U14267 : OAI221_X1 port map( B1 => n1815_port, B2 => n10736, C1 => 
                           n1879_port, C2 => n10727, A => n9242, ZN => n9230);
   U14268 : AOI222_X1 port map( A1 => n10718, A2 => n9688, B1 => n10710, B2 => 
                           n10136, C1 => n10702, C2 => n10584, ZN => n9242);
   U14269 : OAI221_X1 port map( B1 => n1814_port, B2 => n10736, C1 => 
                           n1878_port, C2 => n10727, A => n9260, ZN => n9248);
   U14270 : AOI222_X1 port map( A1 => n10718, A2 => n9689, B1 => n10710, B2 => 
                           n10137, C1 => n10702, C2 => n10585, ZN => n9260);
   U14271 : OAI221_X1 port map( B1 => n1813_port, B2 => n10736, C1 => 
                           n1877_port, C2 => n10727, A => n9278, ZN => n9266);
   U14272 : AOI222_X1 port map( A1 => n10718, A2 => n9690, B1 => n10710, B2 => 
                           n10138, C1 => n10702, C2 => n10586, ZN => n9278);
   U14273 : OAI221_X1 port map( B1 => n1812_port, B2 => n10736, C1 => 
                           n1876_port, C2 => n10727, A => n9296, ZN => n9284);
   U14274 : AOI222_X1 port map( A1 => n10718, A2 => n9691, B1 => n10710, B2 => 
                           n10139, C1 => n10702, C2 => n10587, ZN => n9296);
   U14275 : OAI221_X1 port map( B1 => n1811_port, B2 => n10736, C1 => 
                           n1875_port, C2 => n10727, A => n9314, ZN => n9302);
   U14276 : AOI222_X1 port map( A1 => n10718, A2 => n9692, B1 => n10710, B2 => 
                           n10140, C1 => n10702, C2 => n10588, ZN => n9314);
   U14277 : OAI221_X1 port map( B1 => n1810_port, B2 => n10736, C1 => 
                           n1874_port, C2 => n10727, A => n9332, ZN => n9320);
   U14278 : AOI222_X1 port map( A1 => n10718, A2 => n9693, B1 => n10710, B2 => 
                           n10141, C1 => n10702, C2 => n10589, ZN => n9332);
   U14279 : OAI221_X1 port map( B1 => n1809_port, B2 => n10736, C1 => 
                           n1873_port, C2 => n10727, A => n9350, ZN => n9338);
   U14280 : AOI222_X1 port map( A1 => n10718, A2 => n9694, B1 => n10710, B2 => 
                           n10142, C1 => n10702, C2 => n10590, ZN => n9350);
   U14281 : OAI221_X1 port map( B1 => n1808_port, B2 => n10736, C1 => 
                           n1872_port, C2 => n10727, A => n9368, ZN => n9356);
   U14282 : AOI222_X1 port map( A1 => n10718, A2 => n9695, B1 => n10710, B2 => 
                           n10143, C1 => n10702, C2 => n10591, ZN => n9368);
   U14283 : OAI221_X1 port map( B1 => n1807_port, B2 => n10736, C1 => 
                           n1871_port, C2 => n10727, A => n9386, ZN => n9374);
   U14284 : AOI222_X1 port map( A1 => n10718, A2 => n9696, B1 => n10710, B2 => 
                           n10144, C1 => n10702, C2 => n10592, ZN => n9386);
   U14285 : OAI221_X1 port map( B1 => n1806_port, B2 => n10736, C1 => 
                           n1870_port, C2 => n10727, A => n9404, ZN => n9392);
   U14286 : AOI222_X1 port map( A1 => n10718, A2 => n9697, B1 => n10710, B2 => 
                           n10145, C1 => n10702, C2 => n10593, ZN => n9404);
   U14287 : OAI221_X1 port map( B1 => n1805_port, B2 => n10736, C1 => 
                           n1869_port, C2 => n10727, A => n9422, ZN => n9410);
   U14288 : AOI222_X1 port map( A1 => n10718, A2 => n9698, B1 => n10710, B2 => 
                           n10146, C1 => n10702, C2 => n10594, ZN => n9422);
   U14289 : OAI221_X1 port map( B1 => n1804_port, B2 => n10735, C1 => 
                           n1868_port, C2 => n10726, A => n9440, ZN => n9428);
   U14290 : AOI222_X1 port map( A1 => n10717, A2 => n9699, B1 => n10709, B2 => 
                           n10147, C1 => n10701, C2 => n10595, ZN => n9440);
   U14291 : OAI221_X1 port map( B1 => n1803_port, B2 => n10735, C1 => 
                           n1867_port, C2 => n10726, A => n9458, ZN => n9446);
   U14292 : AOI222_X1 port map( A1 => n10717, A2 => n9700, B1 => n10709, B2 => 
                           n10148, C1 => n10701, C2 => n10596, ZN => n9458);
   U14293 : OAI221_X1 port map( B1 => n1802_port, B2 => n10735, C1 => 
                           n1866_port, C2 => n10726, A => n9476, ZN => n9464);
   U14294 : AOI222_X1 port map( A1 => n10717, A2 => n9701, B1 => n10709, B2 => 
                           n10149, C1 => n10701, C2 => n10597, ZN => n9476);
   U14295 : OAI221_X1 port map( B1 => n1801_port, B2 => n10735, C1 => 
                           n1865_port, C2 => n10726, A => n9494, ZN => n9482);
   U14296 : AOI222_X1 port map( A1 => n10717, A2 => n9702, B1 => n10709, B2 => 
                           n10150, C1 => n10701, C2 => n10598, ZN => n9494);
   U14297 : OAI221_X1 port map( B1 => n1800_port, B2 => n10735, C1 => 
                           n1864_port, C2 => n10726, A => n9512, ZN => n9500);
   U14298 : AOI222_X1 port map( A1 => n10717, A2 => n9703, B1 => n10709, B2 => 
                           n10151, C1 => n10701, C2 => n10599, ZN => n9512);
   U14299 : OAI221_X1 port map( B1 => n1799_port, B2 => n10735, C1 => 
                           n1863_port, C2 => n10726, A => n9530, ZN => n9518);
   U14300 : AOI222_X1 port map( A1 => n10717, A2 => n9704, B1 => n10709, B2 => 
                           n10152, C1 => n10701, C2 => n10600, ZN => n9530);
   U14301 : OAI221_X1 port map( B1 => n1798_port, B2 => n10735, C1 => 
                           n1862_port, C2 => n10726, A => n9548, ZN => n9536);
   U14302 : AOI222_X1 port map( A1 => n10717, A2 => n9705, B1 => n10709, B2 => 
                           n10153, C1 => n10701, C2 => n10601, ZN => n9548);
   U14303 : OAI221_X1 port map( B1 => n1797_port, B2 => n10735, C1 => 
                           n1861_port, C2 => n10726, A => n9566, ZN => n9554);
   U14304 : AOI222_X1 port map( A1 => n10717, A2 => n9706, B1 => n10709, B2 => 
                           n10154, C1 => n10701, C2 => n10602, ZN => n9566);
   U14305 : OAI221_X1 port map( B1 => n1796_port, B2 => n10735, C1 => 
                           n1860_port, C2 => n10726, A => n9584, ZN => n9572);
   U14306 : AOI222_X1 port map( A1 => n10717, A2 => n9707, B1 => n10709, B2 => 
                           n10155, C1 => n10701, C2 => n10603, ZN => n9584);
   U14307 : OAI221_X1 port map( B1 => n1795_port, B2 => n10735, C1 => 
                           n1859_port, C2 => n10726, A => n9602, ZN => n9590);
   U14308 : AOI222_X1 port map( A1 => n10717, A2 => n9708, B1 => n10709, B2 => 
                           n10156, C1 => n10701, C2 => n10604, ZN => n9602);
   U14309 : OAI221_X1 port map( B1 => n1794_port, B2 => n10735, C1 => 
                           n1858_port, C2 => n10726, A => n9620, ZN => n9608);
   U14310 : AOI222_X1 port map( A1 => n10717, A2 => n9709, B1 => n10709, B2 => 
                           n10157, C1 => n10701, C2 => n10605, ZN => n9620);
   U14311 : OAI221_X1 port map( B1 => n1793_port, B2 => n10735, C1 => 
                           n1857_port, C2 => n10726, A => n9643, ZN => n9626);
   U14312 : AOI222_X1 port map( A1 => n10717, A2 => n9710, B1 => n10709, B2 => 
                           n10158, C1 => n10701, C2 => n10606, ZN => n9643);
   U14313 : OAI22_X1 port map( A1 => n320_port, A2 => n11543, B1 => n448_port, 
                           B2 => n11560, ZN => n7299);
   U14314 : OAI22_X1 port map( A1 => n832_port, A2 => n11543, B1 => n960_port, 
                           B2 => n11560, ZN => n7306);
   U14315 : OAI22_X1 port map( A1 => n319_port, A2 => n11543, B1 => n447_port, 
                           B2 => n11560, ZN => n7336);
   U14316 : OAI22_X1 port map( A1 => n831_port, A2 => n11543, B1 => n959_port, 
                           B2 => n11560, ZN => n7340);
   U14317 : OAI22_X1 port map( A1 => n318_port, A2 => n11543, B1 => n446_port, 
                           B2 => n11560, ZN => n7354);
   U14318 : OAI22_X1 port map( A1 => n830_port, A2 => n11543, B1 => n958_port, 
                           B2 => n11560, ZN => n7358);
   U14319 : OAI22_X1 port map( A1 => n317_port, A2 => n11543, B1 => n445_port, 
                           B2 => n11560, ZN => n7372);
   U14320 : OAI22_X1 port map( A1 => n829_port, A2 => n11543, B1 => n957_port, 
                           B2 => n11560, ZN => n7376);
   U14321 : OAI22_X1 port map( A1 => n316_port, A2 => n11542, B1 => n444_port, 
                           B2 => n11559, ZN => n7390);
   U14322 : OAI22_X1 port map( A1 => n828_port, A2 => n11542, B1 => n956_port, 
                           B2 => n11559, ZN => n7394);
   U14323 : OAI22_X1 port map( A1 => n315_port, A2 => n11542, B1 => n443_port, 
                           B2 => n11559, ZN => n7408);
   U14324 : OAI22_X1 port map( A1 => n827_port, A2 => n11542, B1 => n955_port, 
                           B2 => n11559, ZN => n7412);
   U14325 : OAI22_X1 port map( A1 => n314_port, A2 => n11542, B1 => n442_port, 
                           B2 => n11559, ZN => n7426);
   U14326 : OAI22_X1 port map( A1 => n826_port, A2 => n11542, B1 => n954_port, 
                           B2 => n11559, ZN => n7430);
   U14327 : OAI22_X1 port map( A1 => n313_port, A2 => n11542, B1 => n441_port, 
                           B2 => n11559, ZN => n7444);
   U14328 : OAI22_X1 port map( A1 => n825_port, A2 => n11542, B1 => n953_port, 
                           B2 => n11559, ZN => n7448);
   U14329 : OAI22_X1 port map( A1 => n312_port, A2 => n11542, B1 => n440_port, 
                           B2 => n11559, ZN => n7462);
   U14330 : OAI22_X1 port map( A1 => n824_port, A2 => n11542, B1 => n952_port, 
                           B2 => n11559, ZN => n7466);
   U14331 : OAI22_X1 port map( A1 => n311_port, A2 => n11542, B1 => n439_port, 
                           B2 => n11559, ZN => n7480);
   U14332 : OAI22_X1 port map( A1 => n823_port, A2 => n11542, B1 => n951_port, 
                           B2 => n11559, ZN => n7484);
   U14333 : OAI22_X1 port map( A1 => n310_port, A2 => n11541, B1 => n438_port, 
                           B2 => n11558, ZN => n7498);
   U14334 : OAI22_X1 port map( A1 => n822_port, A2 => n11541, B1 => n950_port, 
                           B2 => n11558, ZN => n7502);
   U14335 : OAI22_X1 port map( A1 => n309_port, A2 => n11541, B1 => n437_port, 
                           B2 => n11558, ZN => n7516);
   U14336 : OAI22_X1 port map( A1 => n821_port, A2 => n11541, B1 => n949_port, 
                           B2 => n11558, ZN => n7520);
   U14337 : OAI22_X1 port map( A1 => n308_port, A2 => n11541, B1 => n436_port, 
                           B2 => n11558, ZN => n7534);
   U14338 : OAI22_X1 port map( A1 => n820_port, A2 => n11541, B1 => n948_port, 
                           B2 => n11558, ZN => n7538);
   U14339 : OAI22_X1 port map( A1 => n307_port, A2 => n11541, B1 => n435_port, 
                           B2 => n11558, ZN => n7552);
   U14340 : OAI22_X1 port map( A1 => n819_port, A2 => n11541, B1 => n947_port, 
                           B2 => n11558, ZN => n7556);
   U14341 : OAI22_X1 port map( A1 => n306_port, A2 => n11541, B1 => n434_port, 
                           B2 => n11558, ZN => n7570);
   U14342 : OAI22_X1 port map( A1 => n818_port, A2 => n11541, B1 => n946_port, 
                           B2 => n11558, ZN => n7574);
   U14343 : OAI22_X1 port map( A1 => n305_port, A2 => n11541, B1 => n433_port, 
                           B2 => n11558, ZN => n7588);
   U14344 : OAI22_X1 port map( A1 => n817_port, A2 => n11541, B1 => n945_port, 
                           B2 => n11558, ZN => n7592);
   U14345 : OAI22_X1 port map( A1 => n304_port, A2 => n11540, B1 => n432_port, 
                           B2 => n11557, ZN => n7606);
   U14346 : OAI22_X1 port map( A1 => n816_port, A2 => n11540, B1 => n944_port, 
                           B2 => n11557, ZN => n7610);
   U14347 : OAI22_X1 port map( A1 => n303_port, A2 => n11540, B1 => n431_port, 
                           B2 => n11557, ZN => n7624);
   U14348 : OAI22_X1 port map( A1 => n815_port, A2 => n11540, B1 => n943_port, 
                           B2 => n11557, ZN => n7628);
   U14349 : OAI22_X1 port map( A1 => n302_port, A2 => n11540, B1 => n430_port, 
                           B2 => n11557, ZN => n7642);
   U14350 : OAI22_X1 port map( A1 => n814_port, A2 => n11540, B1 => n942_port, 
                           B2 => n11557, ZN => n7646);
   U14351 : OAI22_X1 port map( A1 => n301_port, A2 => n11540, B1 => n429_port, 
                           B2 => n11557, ZN => n7660);
   U14352 : OAI22_X1 port map( A1 => n813_port, A2 => n11540, B1 => n941_port, 
                           B2 => n11557, ZN => n7664);
   U14353 : OAI22_X1 port map( A1 => n300_port, A2 => n11540, B1 => n428_port, 
                           B2 => n11557, ZN => n7678);
   U14354 : OAI22_X1 port map( A1 => n812_port, A2 => n11540, B1 => n940_port, 
                           B2 => n11557, ZN => n7682);
   U14355 : OAI22_X1 port map( A1 => n299_port, A2 => n11540, B1 => n427_port, 
                           B2 => n11557, ZN => n7696);
   U14356 : OAI22_X1 port map( A1 => n811_port, A2 => n11540, B1 => n939_port, 
                           B2 => n11557, ZN => n7700);
   U14357 : OAI22_X1 port map( A1 => n298_port, A2 => n11539, B1 => n426_port, 
                           B2 => n11556, ZN => n7714);
   U14358 : OAI22_X1 port map( A1 => n810_port, A2 => n11539, B1 => n938_port, 
                           B2 => n11556, ZN => n7718);
   U14359 : OAI22_X1 port map( A1 => n297_port, A2 => n11539, B1 => n425_port, 
                           B2 => n11556, ZN => n7732);
   U14360 : OAI22_X1 port map( A1 => n809_port, A2 => n11539, B1 => n937_port, 
                           B2 => n11556, ZN => n7736);
   U14361 : OAI22_X1 port map( A1 => n296_port, A2 => n11539, B1 => n424_port, 
                           B2 => n11556, ZN => n7750);
   U14362 : OAI22_X1 port map( A1 => n808_port, A2 => n11539, B1 => n936_port, 
                           B2 => n11556, ZN => n7754);
   U14363 : OAI22_X1 port map( A1 => n295_port, A2 => n11539, B1 => n423_port, 
                           B2 => n11556, ZN => n7768);
   U14364 : OAI22_X1 port map( A1 => n807_port, A2 => n11539, B1 => n935_port, 
                           B2 => n11556, ZN => n7772);
   U14365 : OAI22_X1 port map( A1 => n294_port, A2 => n11539, B1 => n422_port, 
                           B2 => n11556, ZN => n7786);
   U14366 : OAI22_X1 port map( A1 => n806_port, A2 => n11539, B1 => n934_port, 
                           B2 => n11556, ZN => n7790);
   U14367 : OAI22_X1 port map( A1 => n293_port, A2 => n11539, B1 => n421_port, 
                           B2 => n11556, ZN => n7804);
   U14368 : OAI22_X1 port map( A1 => n805_port, A2 => n11539, B1 => n933_port, 
                           B2 => n11556, ZN => n7808);
   U14369 : OAI22_X1 port map( A1 => n292_port, A2 => n11538, B1 => n420_port, 
                           B2 => n11555, ZN => n7822);
   U14370 : OAI22_X1 port map( A1 => n804_port, A2 => n11538, B1 => n932_port, 
                           B2 => n11555, ZN => n7826);
   U14371 : OAI22_X1 port map( A1 => n291_port, A2 => n11538, B1 => n419_port, 
                           B2 => n11555, ZN => n7840);
   U14372 : OAI22_X1 port map( A1 => n803_port, A2 => n11538, B1 => n931_port, 
                           B2 => n11555, ZN => n7844);
   U14373 : OAI22_X1 port map( A1 => n290_port, A2 => n11538, B1 => n418_port, 
                           B2 => n11555, ZN => n7858);
   U14374 : OAI22_X1 port map( A1 => n802_port, A2 => n11538, B1 => n930_port, 
                           B2 => n11555, ZN => n7862);
   U14375 : OAI22_X1 port map( A1 => n289_port, A2 => n11538, B1 => n417_port, 
                           B2 => n11555, ZN => n7876);
   U14376 : OAI22_X1 port map( A1 => n801_port, A2 => n11538, B1 => n929_port, 
                           B2 => n11555, ZN => n7880);
   U14377 : OAI22_X1 port map( A1 => n288_port, A2 => n11538, B1 => n416_port, 
                           B2 => n11555, ZN => n7894);
   U14378 : OAI22_X1 port map( A1 => n800_port, A2 => n11538, B1 => n928_port, 
                           B2 => n11555, ZN => n7898);
   U14379 : OAI22_X1 port map( A1 => n287_port, A2 => n11538, B1 => n415_port, 
                           B2 => n11555, ZN => n7912);
   U14380 : OAI22_X1 port map( A1 => n799_port, A2 => n11538, B1 => n927_port, 
                           B2 => n11555, ZN => n7916);
   U14381 : OAI22_X1 port map( A1 => n286_port, A2 => n11537, B1 => n414_port, 
                           B2 => n11554, ZN => n7930);
   U14382 : OAI22_X1 port map( A1 => n798_port, A2 => n11537, B1 => n926_port, 
                           B2 => n11554, ZN => n7934);
   U14383 : OAI22_X1 port map( A1 => n285_port, A2 => n11537, B1 => n413_port, 
                           B2 => n11554, ZN => n7948);
   U14384 : OAI22_X1 port map( A1 => n797_port, A2 => n11537, B1 => n925_port, 
                           B2 => n11554, ZN => n7952);
   U14385 : OAI22_X1 port map( A1 => n284_port, A2 => n11537, B1 => n412_port, 
                           B2 => n11554, ZN => n7966);
   U14386 : OAI22_X1 port map( A1 => n796_port, A2 => n11537, B1 => n924_port, 
                           B2 => n11554, ZN => n7970);
   U14387 : OAI22_X1 port map( A1 => n283_port, A2 => n11537, B1 => n411_port, 
                           B2 => n11554, ZN => n7984);
   U14388 : OAI22_X1 port map( A1 => n795_port, A2 => n11537, B1 => n923_port, 
                           B2 => n11554, ZN => n7988);
   U14389 : OAI22_X1 port map( A1 => n282_port, A2 => n11537, B1 => n410_port, 
                           B2 => n11554, ZN => n8002);
   U14390 : OAI22_X1 port map( A1 => n794_port, A2 => n11537, B1 => n922_port, 
                           B2 => n11554, ZN => n8006);
   U14391 : OAI22_X1 port map( A1 => n281_port, A2 => n11537, B1 => n409_port, 
                           B2 => n11554, ZN => n8020);
   U14392 : OAI22_X1 port map( A1 => n793_port, A2 => n11537, B1 => n921_port, 
                           B2 => n11554, ZN => n8024);
   U14393 : OAI22_X1 port map( A1 => n280_port, A2 => n11536, B1 => n408_port, 
                           B2 => n11553, ZN => n8038);
   U14394 : OAI22_X1 port map( A1 => n792_port, A2 => n11536, B1 => n920_port, 
                           B2 => n11553, ZN => n8042);
   U14395 : OAI22_X1 port map( A1 => n279_port, A2 => n11536, B1 => n407_port, 
                           B2 => n11553, ZN => n8056);
   U14396 : OAI22_X1 port map( A1 => n791_port, A2 => n11536, B1 => n919_port, 
                           B2 => n11553, ZN => n8060);
   U14397 : OAI22_X1 port map( A1 => n278_port, A2 => n11536, B1 => n406_port, 
                           B2 => n11553, ZN => n8074);
   U14398 : OAI22_X1 port map( A1 => n790_port, A2 => n11536, B1 => n918_port, 
                           B2 => n11553, ZN => n8078);
   U14399 : OAI22_X1 port map( A1 => n277_port, A2 => n11536, B1 => n405_port, 
                           B2 => n11553, ZN => n8092);
   U14400 : OAI22_X1 port map( A1 => n789_port, A2 => n11536, B1 => n917_port, 
                           B2 => n11553, ZN => n8096);
   U14401 : OAI22_X1 port map( A1 => n276_port, A2 => n11536, B1 => n404_port, 
                           B2 => n11553, ZN => n8110);
   U14402 : OAI22_X1 port map( A1 => n788_port, A2 => n11536, B1 => n916_port, 
                           B2 => n11553, ZN => n8114);
   U14403 : OAI22_X1 port map( A1 => n275_port, A2 => n11536, B1 => n403_port, 
                           B2 => n11553, ZN => n8128);
   U14404 : OAI22_X1 port map( A1 => n787_port, A2 => n11536, B1 => n915_port, 
                           B2 => n11553, ZN => n8132);
   U14405 : OAI22_X1 port map( A1 => n274_port, A2 => n11535, B1 => n402_port, 
                           B2 => n11552, ZN => n8146);
   U14406 : OAI22_X1 port map( A1 => n786_port, A2 => n11535, B1 => n914_port, 
                           B2 => n11552, ZN => n8150);
   U14407 : OAI22_X1 port map( A1 => n273_port, A2 => n11535, B1 => n401_port, 
                           B2 => n11552, ZN => n8164);
   U14408 : OAI22_X1 port map( A1 => n785_port, A2 => n11535, B1 => n913_port, 
                           B2 => n11552, ZN => n8168);
   U14409 : OAI22_X1 port map( A1 => n272_port, A2 => n11535, B1 => n400_port, 
                           B2 => n11552, ZN => n8182);
   U14410 : OAI22_X1 port map( A1 => n784_port, A2 => n11535, B1 => n912_port, 
                           B2 => n11552, ZN => n8186);
   U14411 : OAI22_X1 port map( A1 => n271_port, A2 => n11535, B1 => n399_port, 
                           B2 => n11552, ZN => n8200);
   U14412 : OAI22_X1 port map( A1 => n783_port, A2 => n11535, B1 => n911_port, 
                           B2 => n11552, ZN => n8204);
   U14413 : OAI22_X1 port map( A1 => n270_port, A2 => n11535, B1 => n398_port, 
                           B2 => n11552, ZN => n8218);
   U14414 : OAI22_X1 port map( A1 => n782_port, A2 => n11535, B1 => n910_port, 
                           B2 => n11552, ZN => n8222);
   U14415 : OAI22_X1 port map( A1 => n269_port, A2 => n11535, B1 => n397_port, 
                           B2 => n11552, ZN => n8236);
   U14416 : OAI22_X1 port map( A1 => n781_port, A2 => n11535, B1 => n909_port, 
                           B2 => n11552, ZN => n8240);
   U14417 : OAI22_X1 port map( A1 => n268_port, A2 => n11534, B1 => n396_port, 
                           B2 => n11551, ZN => n8254);
   U14418 : OAI22_X1 port map( A1 => n780_port, A2 => n11534, B1 => n908_port, 
                           B2 => n11551, ZN => n8258);
   U14419 : OAI22_X1 port map( A1 => n267_port, A2 => n11534, B1 => n395_port, 
                           B2 => n11551, ZN => n8272);
   U14420 : OAI22_X1 port map( A1 => n779_port, A2 => n11534, B1 => n907_port, 
                           B2 => n11551, ZN => n8276);
   U14421 : OAI22_X1 port map( A1 => n266_port, A2 => n11534, B1 => n394_port, 
                           B2 => n11551, ZN => n8290);
   U14422 : OAI22_X1 port map( A1 => n778_port, A2 => n11534, B1 => n906_port, 
                           B2 => n11551, ZN => n8294);
   U14423 : OAI22_X1 port map( A1 => n265_port, A2 => n11534, B1 => n393_port, 
                           B2 => n11551, ZN => n8308);
   U14424 : OAI22_X1 port map( A1 => n777_port, A2 => n11534, B1 => n905_port, 
                           B2 => n11551, ZN => n8312);
   U14425 : OAI22_X1 port map( A1 => n264_port, A2 => n11534, B1 => n392_port, 
                           B2 => n11551, ZN => n8326);
   U14426 : OAI22_X1 port map( A1 => n776_port, A2 => n11534, B1 => n904_port, 
                           B2 => n11551, ZN => n8330);
   U14427 : OAI22_X1 port map( A1 => n263_port, A2 => n11534, B1 => n391_port, 
                           B2 => n11551, ZN => n8344);
   U14428 : OAI22_X1 port map( A1 => n775_port, A2 => n11534, B1 => n903_port, 
                           B2 => n11551, ZN => n8348);
   U14429 : OAI22_X1 port map( A1 => n262_port, A2 => n11533, B1 => n390_port, 
                           B2 => n11550, ZN => n8362);
   U14430 : OAI22_X1 port map( A1 => n774_port, A2 => n11533, B1 => n902_port, 
                           B2 => n11550, ZN => n8366);
   U14431 : OAI22_X1 port map( A1 => n261_port, A2 => n11533, B1 => n389_port, 
                           B2 => n11550, ZN => n8380);
   U14432 : OAI22_X1 port map( A1 => n773_port, A2 => n11533, B1 => n901_port, 
                           B2 => n11550, ZN => n8384);
   U14433 : OAI22_X1 port map( A1 => n260_port, A2 => n11533, B1 => n388_port, 
                           B2 => n11550, ZN => n8398);
   U14434 : OAI22_X1 port map( A1 => n772_port, A2 => n11533, B1 => n900_port, 
                           B2 => n11550, ZN => n8402);
   U14435 : OAI22_X1 port map( A1 => n259_port, A2 => n11533, B1 => n387_port, 
                           B2 => n11550, ZN => n8416);
   U14436 : OAI22_X1 port map( A1 => n771_port, A2 => n11533, B1 => n899_port, 
                           B2 => n11550, ZN => n8420);
   U14437 : OAI22_X1 port map( A1 => n258_port, A2 => n11533, B1 => n386_port, 
                           B2 => n11550, ZN => n8434);
   U14438 : OAI22_X1 port map( A1 => n770_port, A2 => n11533, B1 => n898_port, 
                           B2 => n11550, ZN => n8438);
   U14439 : OAI22_X1 port map( A1 => n257_port, A2 => n11533, B1 => n385_port, 
                           B2 => n11550, ZN => n8452);
   U14440 : OAI22_X1 port map( A1 => n769_port, A2 => n11533, B1 => n897_port, 
                           B2 => n11550, ZN => n8456);
   U14441 : OAI22_X1 port map( A1 => n320_port, A2 => n11611, B1 => n448_port, 
                           B2 => n11628, ZN => n8479);
   U14442 : OAI22_X1 port map( A1 => n832_port, A2 => n11611, B1 => n960_port, 
                           B2 => n11628, ZN => n8486);
   U14443 : OAI22_X1 port map( A1 => n319_port, A2 => n11611, B1 => n447_port, 
                           B2 => n11628, ZN => n8516);
   U14444 : OAI22_X1 port map( A1 => n831_port, A2 => n11611, B1 => n959_port, 
                           B2 => n11628, ZN => n8520);
   U14445 : OAI22_X1 port map( A1 => n318_port, A2 => n11611, B1 => n446_port, 
                           B2 => n11628, ZN => n8534);
   U14446 : OAI22_X1 port map( A1 => n830_port, A2 => n11611, B1 => n958_port, 
                           B2 => n11628, ZN => n8538);
   U14447 : OAI22_X1 port map( A1 => n317_port, A2 => n11611, B1 => n445_port, 
                           B2 => n11628, ZN => n8552);
   U14448 : OAI22_X1 port map( A1 => n829_port, A2 => n11611, B1 => n957_port, 
                           B2 => n11628, ZN => n8556);
   U14449 : OAI22_X1 port map( A1 => n316_port, A2 => n11610, B1 => n444_port, 
                           B2 => n11627, ZN => n8570);
   U14450 : OAI22_X1 port map( A1 => n828_port, A2 => n11610, B1 => n956_port, 
                           B2 => n11627, ZN => n8574);
   U14451 : OAI22_X1 port map( A1 => n315_port, A2 => n11610, B1 => n443_port, 
                           B2 => n11627, ZN => n8588);
   U14452 : OAI22_X1 port map( A1 => n827_port, A2 => n11610, B1 => n955_port, 
                           B2 => n11627, ZN => n8592);
   U14453 : OAI22_X1 port map( A1 => n314_port, A2 => n11610, B1 => n442_port, 
                           B2 => n11627, ZN => n8606);
   U14454 : OAI22_X1 port map( A1 => n826_port, A2 => n11610, B1 => n954_port, 
                           B2 => n11627, ZN => n8610);
   U14455 : OAI22_X1 port map( A1 => n313_port, A2 => n11610, B1 => n441_port, 
                           B2 => n11627, ZN => n8624);
   U14456 : OAI22_X1 port map( A1 => n825_port, A2 => n11610, B1 => n953_port, 
                           B2 => n11627, ZN => n8628);
   U14457 : OAI22_X1 port map( A1 => n312_port, A2 => n11610, B1 => n440_port, 
                           B2 => n11627, ZN => n8642);
   U14458 : OAI22_X1 port map( A1 => n824_port, A2 => n11610, B1 => n952_port, 
                           B2 => n11627, ZN => n8646);
   U14459 : OAI22_X1 port map( A1 => n311_port, A2 => n11610, B1 => n439_port, 
                           B2 => n11627, ZN => n8660);
   U14460 : OAI22_X1 port map( A1 => n823_port, A2 => n11610, B1 => n951_port, 
                           B2 => n11627, ZN => n8664);
   U14461 : OAI22_X1 port map( A1 => n310_port, A2 => n11609, B1 => n438_port, 
                           B2 => n11626, ZN => n8678);
   U14462 : OAI22_X1 port map( A1 => n822_port, A2 => n11609, B1 => n950_port, 
                           B2 => n11626, ZN => n8682);
   U14463 : OAI22_X1 port map( A1 => n309_port, A2 => n11609, B1 => n437_port, 
                           B2 => n11626, ZN => n8696);
   U14464 : OAI22_X1 port map( A1 => n821_port, A2 => n11609, B1 => n949_port, 
                           B2 => n11626, ZN => n8700);
   U14465 : OAI22_X1 port map( A1 => n308_port, A2 => n11609, B1 => n436_port, 
                           B2 => n11626, ZN => n8714);
   U14466 : OAI22_X1 port map( A1 => n820_port, A2 => n11609, B1 => n948_port, 
                           B2 => n11626, ZN => n8718);
   U14467 : OAI22_X1 port map( A1 => n307_port, A2 => n11609, B1 => n435_port, 
                           B2 => n11626, ZN => n8732);
   U14468 : OAI22_X1 port map( A1 => n819_port, A2 => n11609, B1 => n947_port, 
                           B2 => n11626, ZN => n8736);
   U14469 : OAI22_X1 port map( A1 => n306_port, A2 => n11609, B1 => n434_port, 
                           B2 => n11626, ZN => n8750);
   U14470 : OAI22_X1 port map( A1 => n818_port, A2 => n11609, B1 => n946_port, 
                           B2 => n11626, ZN => n8754);
   U14471 : OAI22_X1 port map( A1 => n305_port, A2 => n11609, B1 => n433_port, 
                           B2 => n11626, ZN => n8768);
   U14472 : OAI22_X1 port map( A1 => n817_port, A2 => n11609, B1 => n945_port, 
                           B2 => n11626, ZN => n8772);
   U14473 : OAI22_X1 port map( A1 => n304_port, A2 => n11608, B1 => n432_port, 
                           B2 => n11625, ZN => n8786);
   U14474 : OAI22_X1 port map( A1 => n816_port, A2 => n11608, B1 => n944_port, 
                           B2 => n11625, ZN => n8790);
   U14475 : OAI22_X1 port map( A1 => n303_port, A2 => n11608, B1 => n431_port, 
                           B2 => n11625, ZN => n8804);
   U14476 : OAI22_X1 port map( A1 => n815_port, A2 => n11608, B1 => n943_port, 
                           B2 => n11625, ZN => n8808);
   U14477 : OAI22_X1 port map( A1 => n302_port, A2 => n11608, B1 => n430_port, 
                           B2 => n11625, ZN => n8822);
   U14478 : OAI22_X1 port map( A1 => n814_port, A2 => n11608, B1 => n942_port, 
                           B2 => n11625, ZN => n8826);
   U14479 : OAI22_X1 port map( A1 => n301_port, A2 => n11608, B1 => n429_port, 
                           B2 => n11625, ZN => n8840);
   U14480 : OAI22_X1 port map( A1 => n813_port, A2 => n11608, B1 => n941_port, 
                           B2 => n11625, ZN => n8844);
   U14481 : OAI22_X1 port map( A1 => n300_port, A2 => n11608, B1 => n428_port, 
                           B2 => n11625, ZN => n8858);
   U14482 : OAI22_X1 port map( A1 => n812_port, A2 => n11608, B1 => n940_port, 
                           B2 => n11625, ZN => n8862);
   U14483 : OAI22_X1 port map( A1 => n299_port, A2 => n11608, B1 => n427_port, 
                           B2 => n11625, ZN => n8876);
   U14484 : OAI22_X1 port map( A1 => n811_port, A2 => n11608, B1 => n939_port, 
                           B2 => n11625, ZN => n8880);
   U14485 : OAI22_X1 port map( A1 => n298_port, A2 => n11607, B1 => n426_port, 
                           B2 => n11624, ZN => n8894);
   U14486 : OAI22_X1 port map( A1 => n810_port, A2 => n11607, B1 => n938_port, 
                           B2 => n11624, ZN => n8898);
   U14487 : OAI22_X1 port map( A1 => n297_port, A2 => n11607, B1 => n425_port, 
                           B2 => n11624, ZN => n8912);
   U14488 : OAI22_X1 port map( A1 => n809_port, A2 => n11607, B1 => n937_port, 
                           B2 => n11624, ZN => n8916);
   U14489 : OAI22_X1 port map( A1 => n296_port, A2 => n11607, B1 => n424_port, 
                           B2 => n11624, ZN => n8930);
   U14490 : OAI22_X1 port map( A1 => n808_port, A2 => n11607, B1 => n936_port, 
                           B2 => n11624, ZN => n8934);
   U14491 : OAI22_X1 port map( A1 => n295_port, A2 => n11607, B1 => n423_port, 
                           B2 => n11624, ZN => n8948);
   U14492 : OAI22_X1 port map( A1 => n807_port, A2 => n11607, B1 => n935_port, 
                           B2 => n11624, ZN => n8952);
   U14493 : OAI22_X1 port map( A1 => n294_port, A2 => n11607, B1 => n422_port, 
                           B2 => n11624, ZN => n8966);
   U14494 : OAI22_X1 port map( A1 => n806_port, A2 => n11607, B1 => n934_port, 
                           B2 => n11624, ZN => n8970);
   U14495 : OAI22_X1 port map( A1 => n293_port, A2 => n11607, B1 => n421_port, 
                           B2 => n11624, ZN => n8984);
   U14496 : OAI22_X1 port map( A1 => n805_port, A2 => n11607, B1 => n933_port, 
                           B2 => n11624, ZN => n8988);
   U14497 : OAI22_X1 port map( A1 => n292_port, A2 => n11606, B1 => n420_port, 
                           B2 => n11623, ZN => n9002);
   U14498 : OAI22_X1 port map( A1 => n804_port, A2 => n11606, B1 => n932_port, 
                           B2 => n11623, ZN => n9006);
   U14499 : OAI22_X1 port map( A1 => n291_port, A2 => n11606, B1 => n419_port, 
                           B2 => n11623, ZN => n9020);
   U14500 : OAI22_X1 port map( A1 => n803_port, A2 => n11606, B1 => n931_port, 
                           B2 => n11623, ZN => n9024);
   U14501 : OAI22_X1 port map( A1 => n290_port, A2 => n11606, B1 => n418_port, 
                           B2 => n11623, ZN => n9038);
   U14502 : OAI22_X1 port map( A1 => n802_port, A2 => n11606, B1 => n930_port, 
                           B2 => n11623, ZN => n9042);
   U14503 : OAI22_X1 port map( A1 => n289_port, A2 => n11606, B1 => n417_port, 
                           B2 => n11623, ZN => n9056);
   U14504 : OAI22_X1 port map( A1 => n801_port, A2 => n11606, B1 => n929_port, 
                           B2 => n11623, ZN => n9060);
   U14505 : OAI22_X1 port map( A1 => n288_port, A2 => n11606, B1 => n416_port, 
                           B2 => n11623, ZN => n9074);
   U14506 : OAI22_X1 port map( A1 => n800_port, A2 => n11606, B1 => n928_port, 
                           B2 => n11623, ZN => n9078);
   U14507 : OAI22_X1 port map( A1 => n287_port, A2 => n11606, B1 => n415_port, 
                           B2 => n11623, ZN => n9092);
   U14508 : OAI22_X1 port map( A1 => n799_port, A2 => n11606, B1 => n927_port, 
                           B2 => n11623, ZN => n9096);
   U14509 : OAI22_X1 port map( A1 => n286_port, A2 => n11605, B1 => n414_port, 
                           B2 => n11622, ZN => n9110);
   U14510 : OAI22_X1 port map( A1 => n798_port, A2 => n11605, B1 => n926_port, 
                           B2 => n11622, ZN => n9114);
   U14511 : OAI22_X1 port map( A1 => n285_port, A2 => n11605, B1 => n413_port, 
                           B2 => n11622, ZN => n9128);
   U14512 : OAI22_X1 port map( A1 => n797_port, A2 => n11605, B1 => n925_port, 
                           B2 => n11622, ZN => n9132);
   U14513 : OAI22_X1 port map( A1 => n284_port, A2 => n11605, B1 => n412_port, 
                           B2 => n11622, ZN => n9146);
   U14514 : OAI22_X1 port map( A1 => n796_port, A2 => n11605, B1 => n924_port, 
                           B2 => n11622, ZN => n9150);
   U14515 : OAI22_X1 port map( A1 => n283_port, A2 => n11605, B1 => n411_port, 
                           B2 => n11622, ZN => n9164);
   U14516 : OAI22_X1 port map( A1 => n795_port, A2 => n11605, B1 => n923_port, 
                           B2 => n11622, ZN => n9168);
   U14517 : OAI22_X1 port map( A1 => n282_port, A2 => n11605, B1 => n410_port, 
                           B2 => n11622, ZN => n9182);
   U14518 : OAI22_X1 port map( A1 => n794_port, A2 => n11605, B1 => n922_port, 
                           B2 => n11622, ZN => n9186);
   U14519 : OAI22_X1 port map( A1 => n281_port, A2 => n11605, B1 => n409_port, 
                           B2 => n11622, ZN => n9200);
   U14520 : OAI22_X1 port map( A1 => n793_port, A2 => n11605, B1 => n921_port, 
                           B2 => n11622, ZN => n9204);
   U14521 : OAI22_X1 port map( A1 => n280_port, A2 => n11604, B1 => n408_port, 
                           B2 => n11621, ZN => n9218);
   U14522 : OAI22_X1 port map( A1 => n792_port, A2 => n11604, B1 => n920_port, 
                           B2 => n11621, ZN => n9222);
   U14523 : OAI22_X1 port map( A1 => n279_port, A2 => n11604, B1 => n407_port, 
                           B2 => n11621, ZN => n9236);
   U14524 : OAI22_X1 port map( A1 => n791_port, A2 => n11604, B1 => n919_port, 
                           B2 => n11621, ZN => n9240);
   U14525 : OAI22_X1 port map( A1 => n278_port, A2 => n11604, B1 => n406_port, 
                           B2 => n11621, ZN => n9254);
   U14526 : OAI22_X1 port map( A1 => n790_port, A2 => n11604, B1 => n918_port, 
                           B2 => n11621, ZN => n9258);
   U14527 : OAI22_X1 port map( A1 => n277_port, A2 => n11604, B1 => n405_port, 
                           B2 => n11621, ZN => n9272);
   U14528 : OAI22_X1 port map( A1 => n789_port, A2 => n11604, B1 => n917_port, 
                           B2 => n11621, ZN => n9276);
   U14529 : OAI22_X1 port map( A1 => n276_port, A2 => n11604, B1 => n404_port, 
                           B2 => n11621, ZN => n9290);
   U14530 : OAI22_X1 port map( A1 => n788_port, A2 => n11604, B1 => n916_port, 
                           B2 => n11621, ZN => n9294);
   U14531 : OAI22_X1 port map( A1 => n275_port, A2 => n11604, B1 => n403_port, 
                           B2 => n11621, ZN => n9308);
   U14532 : OAI22_X1 port map( A1 => n787_port, A2 => n11604, B1 => n915_port, 
                           B2 => n11621, ZN => n9312);
   U14533 : OAI22_X1 port map( A1 => n274_port, A2 => n11603, B1 => n402_port, 
                           B2 => n11620, ZN => n9326);
   U14534 : OAI22_X1 port map( A1 => n786_port, A2 => n11603, B1 => n914_port, 
                           B2 => n11620, ZN => n9330);
   U14535 : OAI22_X1 port map( A1 => n273_port, A2 => n11603, B1 => n401_port, 
                           B2 => n11620, ZN => n9344);
   U14536 : OAI22_X1 port map( A1 => n785_port, A2 => n11603, B1 => n913_port, 
                           B2 => n11620, ZN => n9348);
   U14537 : OAI22_X1 port map( A1 => n272_port, A2 => n11603, B1 => n400_port, 
                           B2 => n11620, ZN => n9362);
   U14538 : OAI22_X1 port map( A1 => n784_port, A2 => n11603, B1 => n912_port, 
                           B2 => n11620, ZN => n9366);
   U14539 : OAI22_X1 port map( A1 => n271_port, A2 => n11603, B1 => n399_port, 
                           B2 => n11620, ZN => n9380);
   U14540 : OAI22_X1 port map( A1 => n783_port, A2 => n11603, B1 => n911_port, 
                           B2 => n11620, ZN => n9384);
   U14541 : OAI22_X1 port map( A1 => n270_port, A2 => n11603, B1 => n398_port, 
                           B2 => n11620, ZN => n9398);
   U14542 : OAI22_X1 port map( A1 => n782_port, A2 => n11603, B1 => n910_port, 
                           B2 => n11620, ZN => n9402);
   U14543 : OAI22_X1 port map( A1 => n269_port, A2 => n11603, B1 => n397_port, 
                           B2 => n11620, ZN => n9416);
   U14544 : OAI22_X1 port map( A1 => n781_port, A2 => n11603, B1 => n909_port, 
                           B2 => n11620, ZN => n9420);
   U14545 : OAI22_X1 port map( A1 => n268_port, A2 => n11602, B1 => n396_port, 
                           B2 => n11619, ZN => n9434);
   U14546 : OAI22_X1 port map( A1 => n780_port, A2 => n11602, B1 => n908_port, 
                           B2 => n11619, ZN => n9438);
   U14547 : OAI22_X1 port map( A1 => n267_port, A2 => n11602, B1 => n395_port, 
                           B2 => n11619, ZN => n9452);
   U14548 : OAI22_X1 port map( A1 => n779_port, A2 => n11602, B1 => n907_port, 
                           B2 => n11619, ZN => n9456);
   U14549 : OAI22_X1 port map( A1 => n266_port, A2 => n11602, B1 => n394_port, 
                           B2 => n11619, ZN => n9470);
   U14550 : OAI22_X1 port map( A1 => n778_port, A2 => n11602, B1 => n906_port, 
                           B2 => n11619, ZN => n9474);
   U14551 : OAI22_X1 port map( A1 => n265_port, A2 => n11602, B1 => n393_port, 
                           B2 => n11619, ZN => n9488);
   U14552 : OAI22_X1 port map( A1 => n777_port, A2 => n11602, B1 => n905_port, 
                           B2 => n11619, ZN => n9492);
   U14553 : OAI22_X1 port map( A1 => n264_port, A2 => n11602, B1 => n392_port, 
                           B2 => n11619, ZN => n9506);
   U14554 : OAI22_X1 port map( A1 => n776_port, A2 => n11602, B1 => n904_port, 
                           B2 => n11619, ZN => n9510);
   U14555 : OAI22_X1 port map( A1 => n263_port, A2 => n11602, B1 => n391_port, 
                           B2 => n11619, ZN => n9524);
   U14556 : OAI22_X1 port map( A1 => n775_port, A2 => n11602, B1 => n903_port, 
                           B2 => n11619, ZN => n9528);
   U14557 : OAI22_X1 port map( A1 => n262_port, A2 => n11601, B1 => n390_port, 
                           B2 => n11618, ZN => n9542);
   U14558 : OAI22_X1 port map( A1 => n774_port, A2 => n11601, B1 => n902_port, 
                           B2 => n11618, ZN => n9546);
   U14559 : OAI22_X1 port map( A1 => n261_port, A2 => n11601, B1 => n389_port, 
                           B2 => n11618, ZN => n9560);
   U14560 : OAI22_X1 port map( A1 => n773_port, A2 => n11601, B1 => n901_port, 
                           B2 => n11618, ZN => n9564);
   U14561 : OAI22_X1 port map( A1 => n260_port, A2 => n11601, B1 => n388_port, 
                           B2 => n11618, ZN => n9578);
   U14562 : OAI22_X1 port map( A1 => n772_port, A2 => n11601, B1 => n900_port, 
                           B2 => n11618, ZN => n9582);
   U14563 : OAI22_X1 port map( A1 => n259_port, A2 => n11601, B1 => n387_port, 
                           B2 => n11618, ZN => n9596);
   U14564 : OAI22_X1 port map( A1 => n771_port, A2 => n11601, B1 => n899_port, 
                           B2 => n11618, ZN => n9600);
   U14565 : OAI22_X1 port map( A1 => n258_port, A2 => n11601, B1 => n386_port, 
                           B2 => n11618, ZN => n9614);
   U14566 : OAI22_X1 port map( A1 => n770_port, A2 => n11601, B1 => n898_port, 
                           B2 => n11618, ZN => n9618);
   U14567 : OAI22_X1 port map( A1 => n257_port, A2 => n11601, B1 => n385_port, 
                           B2 => n11618, ZN => n9632);
   U14568 : OAI22_X1 port map( A1 => n769_port, A2 => n11601, B1 => n897_port, 
                           B2 => n11618, ZN => n9636);
   U14569 : OAI22_X1 port map( A1 => n1472_port, A2 => n10864, B1 => n1408_port
                           , B2 => n10855, ZN => n7324);
   U14570 : OAI22_X1 port map( A1 => n1471_port, A2 => n10864, B1 => n1407_port
                           , B2 => n10855, ZN => n7344);
   U14571 : OAI22_X1 port map( A1 => n1470_port, A2 => n10864, B1 => n1406_port
                           , B2 => n10855, ZN => n7362);
   U14572 : OAI22_X1 port map( A1 => n1469_port, A2 => n10864, B1 => n1405_port
                           , B2 => n10855, ZN => n7380);
   U14573 : OAI22_X1 port map( A1 => n1468_port, A2 => n10863, B1 => n1404_port
                           , B2 => n10854, ZN => n7398);
   U14574 : OAI22_X1 port map( A1 => n1467_port, A2 => n10863, B1 => n1403_port
                           , B2 => n10854, ZN => n7416);
   U14575 : OAI22_X1 port map( A1 => n1466_port, A2 => n10863, B1 => n1402_port
                           , B2 => n10854, ZN => n7434);
   U14576 : OAI22_X1 port map( A1 => n1465_port, A2 => n10863, B1 => n1401_port
                           , B2 => n10854, ZN => n7452);
   U14577 : OAI22_X1 port map( A1 => n1464_port, A2 => n10863, B1 => n1400_port
                           , B2 => n10854, ZN => n7470);
   U14578 : OAI22_X1 port map( A1 => n1463_port, A2 => n10863, B1 => n1399_port
                           , B2 => n10854, ZN => n7488);
   U14579 : OAI22_X1 port map( A1 => n1462_port, A2 => n10863, B1 => n1398_port
                           , B2 => n10854, ZN => n7506);
   U14580 : OAI22_X1 port map( A1 => n1461_port, A2 => n10863, B1 => n1397_port
                           , B2 => n10854, ZN => n7524);
   U14581 : OAI22_X1 port map( A1 => n1460_port, A2 => n10863, B1 => n1396_port
                           , B2 => n10854, ZN => n7542);
   U14582 : OAI22_X1 port map( A1 => n1459_port, A2 => n10863, B1 => n1395_port
                           , B2 => n10854, ZN => n7560);
   U14583 : OAI22_X1 port map( A1 => n1458_port, A2 => n10863, B1 => n1394_port
                           , B2 => n10854, ZN => n7578);
   U14584 : OAI22_X1 port map( A1 => n1457_port, A2 => n10863, B1 => n1393_port
                           , B2 => n10854, ZN => n7596);
   U14585 : OAI22_X1 port map( A1 => n1456_port, A2 => n10862, B1 => n1392_port
                           , B2 => n10853, ZN => n7614);
   U14586 : OAI22_X1 port map( A1 => n1455_port, A2 => n10862, B1 => n1391_port
                           , B2 => n10853, ZN => n7632);
   U14587 : OAI22_X1 port map( A1 => n1454_port, A2 => n10862, B1 => n1390_port
                           , B2 => n10853, ZN => n7650);
   U14588 : OAI22_X1 port map( A1 => n1453_port, A2 => n10862, B1 => n1389_port
                           , B2 => n10853, ZN => n7668);
   U14589 : OAI22_X1 port map( A1 => n1452_port, A2 => n10862, B1 => n1388_port
                           , B2 => n10853, ZN => n7686);
   U14590 : OAI22_X1 port map( A1 => n1451_port, A2 => n10862, B1 => n1387_port
                           , B2 => n10853, ZN => n7704);
   U14591 : OAI22_X1 port map( A1 => n1450_port, A2 => n10862, B1 => n1386_port
                           , B2 => n10853, ZN => n7722);
   U14592 : OAI22_X1 port map( A1 => n1449_port, A2 => n10862, B1 => n1385_port
                           , B2 => n10853, ZN => n7740);
   U14593 : OAI22_X1 port map( A1 => n1448_port, A2 => n10862, B1 => n1384_port
                           , B2 => n10853, ZN => n7758);
   U14594 : OAI22_X1 port map( A1 => n1447_port, A2 => n10862, B1 => n1383_port
                           , B2 => n10853, ZN => n7776);
   U14595 : OAI22_X1 port map( A1 => n1446_port, A2 => n10862, B1 => n1382_port
                           , B2 => n10853, ZN => n7794);
   U14596 : OAI22_X1 port map( A1 => n1445_port, A2 => n10862, B1 => n1381_port
                           , B2 => n10853, ZN => n7812);
   U14597 : OAI22_X1 port map( A1 => n1444_port, A2 => n10861, B1 => n1380_port
                           , B2 => n10852, ZN => n7830);
   U14598 : OAI22_X1 port map( A1 => n1443_port, A2 => n10861, B1 => n1379_port
                           , B2 => n10852, ZN => n7848);
   U14599 : OAI22_X1 port map( A1 => n1442_port, A2 => n10861, B1 => n1378_port
                           , B2 => n10852, ZN => n7866);
   U14600 : OAI22_X1 port map( A1 => n1441_port, A2 => n10861, B1 => n1377_port
                           , B2 => n10852, ZN => n7884);
   U14601 : OAI22_X1 port map( A1 => n1440_port, A2 => n10861, B1 => n1376_port
                           , B2 => n10852, ZN => n7902);
   U14602 : OAI22_X1 port map( A1 => n1439_port, A2 => n10861, B1 => n1375_port
                           , B2 => n10852, ZN => n7920);
   U14603 : OAI22_X1 port map( A1 => n1438_port, A2 => n10861, B1 => n1374_port
                           , B2 => n10852, ZN => n7938);
   U14604 : OAI22_X1 port map( A1 => n1437_port, A2 => n10861, B1 => n1373_port
                           , B2 => n10852, ZN => n7956);
   U14605 : OAI22_X1 port map( A1 => n1436_port, A2 => n10861, B1 => n1372_port
                           , B2 => n10852, ZN => n7974);
   U14606 : OAI22_X1 port map( A1 => n1435_port, A2 => n10861, B1 => n1371_port
                           , B2 => n10852, ZN => n7992);
   U14607 : OAI22_X1 port map( A1 => n1434_port, A2 => n10861, B1 => n1370_port
                           , B2 => n10852, ZN => n8010);
   U14608 : OAI22_X1 port map( A1 => n1433_port, A2 => n10861, B1 => n1369_port
                           , B2 => n10852, ZN => n8028);
   U14609 : OAI22_X1 port map( A1 => n1432_port, A2 => n10860, B1 => n1368_port
                           , B2 => n10851, ZN => n8046);
   U14610 : OAI22_X1 port map( A1 => n1431_port, A2 => n10860, B1 => n1367_port
                           , B2 => n10851, ZN => n8064);
   U14611 : OAI22_X1 port map( A1 => n1430_port, A2 => n10860, B1 => n1366_port
                           , B2 => n10851, ZN => n8082);
   U14612 : OAI22_X1 port map( A1 => n1429_port, A2 => n10860, B1 => n1365_port
                           , B2 => n10851, ZN => n8100);
   U14613 : OAI22_X1 port map( A1 => n1428_port, A2 => n10860, B1 => n1364_port
                           , B2 => n10851, ZN => n8118);
   U14614 : OAI22_X1 port map( A1 => n1427_port, A2 => n10860, B1 => n1363_port
                           , B2 => n10851, ZN => n8136);
   U14615 : OAI22_X1 port map( A1 => n1426_port, A2 => n10860, B1 => n1362_port
                           , B2 => n10851, ZN => n8154);
   U14616 : OAI22_X1 port map( A1 => n1425_port, A2 => n10860, B1 => n1361_port
                           , B2 => n10851, ZN => n8172);
   U14617 : OAI22_X1 port map( A1 => n1424_port, A2 => n10860, B1 => n1360_port
                           , B2 => n10851, ZN => n8190);
   U14618 : OAI22_X1 port map( A1 => n1423_port, A2 => n10860, B1 => n1359_port
                           , B2 => n10851, ZN => n8208);
   U14619 : OAI22_X1 port map( A1 => n1422_port, A2 => n10860, B1 => n1358_port
                           , B2 => n10851, ZN => n8226);
   U14620 : OAI22_X1 port map( A1 => n1421_port, A2 => n10860, B1 => n1357_port
                           , B2 => n10851, ZN => n8244);
   U14621 : OAI22_X1 port map( A1 => n1420_port, A2 => n10859, B1 => n1356_port
                           , B2 => n10850, ZN => n8262);
   U14622 : OAI22_X1 port map( A1 => n1419_port, A2 => n10859, B1 => n1355_port
                           , B2 => n10850, ZN => n8280);
   U14623 : OAI22_X1 port map( A1 => n1418_port, A2 => n10859, B1 => n1354_port
                           , B2 => n10850, ZN => n8298);
   U14624 : OAI22_X1 port map( A1 => n1417_port, A2 => n10859, B1 => n1353_port
                           , B2 => n10850, ZN => n8316);
   U14625 : OAI22_X1 port map( A1 => n1416_port, A2 => n10859, B1 => n1352_port
                           , B2 => n10850, ZN => n8334);
   U14626 : OAI22_X1 port map( A1 => n1415_port, A2 => n10859, B1 => n1351_port
                           , B2 => n10850, ZN => n8352);
   U14627 : OAI22_X1 port map( A1 => n1414_port, A2 => n10859, B1 => n1350_port
                           , B2 => n10850, ZN => n8370);
   U14628 : OAI22_X1 port map( A1 => n1413_port, A2 => n10859, B1 => n1349_port
                           , B2 => n10850, ZN => n8388);
   U14629 : OAI22_X1 port map( A1 => n1412_port, A2 => n10859, B1 => n1348_port
                           , B2 => n10850, ZN => n8406);
   U14630 : OAI22_X1 port map( A1 => n1411_port, A2 => n10859, B1 => n1347_port
                           , B2 => n10850, ZN => n8424);
   U14631 : OAI22_X1 port map( A1 => n1410_port, A2 => n10859, B1 => n1346_port
                           , B2 => n10850, ZN => n8442);
   U14632 : OAI22_X1 port map( A1 => n1409_port, A2 => n10859, B1 => n1345_port
                           , B2 => n10850, ZN => n8466);
   U14633 : OAI22_X1 port map( A1 => n1472_port, A2 => n10639, B1 => n1408_port
                           , B2 => n10630, ZN => n8504);
   U14634 : OAI22_X1 port map( A1 => n1471_port, A2 => n10639, B1 => n1407_port
                           , B2 => n10630, ZN => n8524);
   U14635 : OAI22_X1 port map( A1 => n1470_port, A2 => n10639, B1 => n1406_port
                           , B2 => n10630, ZN => n8542);
   U14636 : OAI22_X1 port map( A1 => n1469_port, A2 => n10639, B1 => n1405_port
                           , B2 => n10630, ZN => n8560);
   U14637 : OAI22_X1 port map( A1 => n1468_port, A2 => n10638, B1 => n1404_port
                           , B2 => n10629, ZN => n8578);
   U14638 : OAI22_X1 port map( A1 => n1467_port, A2 => n10638, B1 => n1403_port
                           , B2 => n10629, ZN => n8596);
   U14639 : OAI22_X1 port map( A1 => n1466_port, A2 => n10638, B1 => n1402_port
                           , B2 => n10629, ZN => n8614);
   U14640 : OAI22_X1 port map( A1 => n1465_port, A2 => n10638, B1 => n1401_port
                           , B2 => n10629, ZN => n8632);
   U14641 : OAI22_X1 port map( A1 => n1464_port, A2 => n10638, B1 => n1400_port
                           , B2 => n10629, ZN => n8650);
   U14642 : OAI22_X1 port map( A1 => n1463_port, A2 => n10638, B1 => n1399_port
                           , B2 => n10629, ZN => n8668);
   U14643 : OAI22_X1 port map( A1 => n1462_port, A2 => n10638, B1 => n1398_port
                           , B2 => n10629, ZN => n8686);
   U14644 : OAI22_X1 port map( A1 => n1461_port, A2 => n10638, B1 => n1397_port
                           , B2 => n10629, ZN => n8704);
   U14645 : OAI22_X1 port map( A1 => n1460_port, A2 => n10638, B1 => n1396_port
                           , B2 => n10629, ZN => n8722);
   U14646 : OAI22_X1 port map( A1 => n1459_port, A2 => n10638, B1 => n1395_port
                           , B2 => n10629, ZN => n8740);
   U14647 : OAI22_X1 port map( A1 => n1458_port, A2 => n10638, B1 => n1394_port
                           , B2 => n10629, ZN => n8758);
   U14648 : OAI22_X1 port map( A1 => n1457_port, A2 => n10638, B1 => n1393_port
                           , B2 => n10629, ZN => n8776);
   U14649 : OAI22_X1 port map( A1 => n1456_port, A2 => n10637, B1 => n1392_port
                           , B2 => n10628, ZN => n8794);
   U14650 : OAI22_X1 port map( A1 => n1455_port, A2 => n10637, B1 => n1391_port
                           , B2 => n10628, ZN => n8812);
   U14651 : OAI22_X1 port map( A1 => n1454_port, A2 => n10637, B1 => n1390_port
                           , B2 => n10628, ZN => n8830);
   U14652 : OAI22_X1 port map( A1 => n1453_port, A2 => n10637, B1 => n1389_port
                           , B2 => n10628, ZN => n8848);
   U14653 : OAI22_X1 port map( A1 => n1452_port, A2 => n10637, B1 => n1388_port
                           , B2 => n10628, ZN => n8866);
   U14654 : OAI22_X1 port map( A1 => n1451_port, A2 => n10637, B1 => n1387_port
                           , B2 => n10628, ZN => n8884);
   U14655 : OAI22_X1 port map( A1 => n1450_port, A2 => n10637, B1 => n1386_port
                           , B2 => n10628, ZN => n8902);
   U14656 : OAI22_X1 port map( A1 => n1449_port, A2 => n10637, B1 => n1385_port
                           , B2 => n10628, ZN => n8920);
   U14657 : OAI22_X1 port map( A1 => n1448_port, A2 => n10637, B1 => n1384_port
                           , B2 => n10628, ZN => n8938);
   U14658 : OAI22_X1 port map( A1 => n1447_port, A2 => n10637, B1 => n1383_port
                           , B2 => n10628, ZN => n8956);
   U14659 : OAI22_X1 port map( A1 => n1446_port, A2 => n10637, B1 => n1382_port
                           , B2 => n10628, ZN => n8974);
   U14660 : OAI22_X1 port map( A1 => n1445_port, A2 => n10637, B1 => n1381_port
                           , B2 => n10628, ZN => n8992);
   U14661 : OAI22_X1 port map( A1 => n1444_port, A2 => n10636, B1 => n1380_port
                           , B2 => n10627, ZN => n9010);
   U14662 : OAI22_X1 port map( A1 => n1443_port, A2 => n10636, B1 => n1379_port
                           , B2 => n10627, ZN => n9028);
   U14663 : OAI22_X1 port map( A1 => n1442_port, A2 => n10636, B1 => n1378_port
                           , B2 => n10627, ZN => n9046);
   U14664 : OAI22_X1 port map( A1 => n1441_port, A2 => n10636, B1 => n1377_port
                           , B2 => n10627, ZN => n9064);
   U14665 : OAI22_X1 port map( A1 => n1440_port, A2 => n10636, B1 => n1376_port
                           , B2 => n10627, ZN => n9082);
   U14666 : OAI22_X1 port map( A1 => n1439_port, A2 => n10636, B1 => n1375_port
                           , B2 => n10627, ZN => n9100);
   U14667 : OAI22_X1 port map( A1 => n1438_port, A2 => n10636, B1 => n1374_port
                           , B2 => n10627, ZN => n9118);
   U14668 : OAI22_X1 port map( A1 => n1437_port, A2 => n10636, B1 => n1373_port
                           , B2 => n10627, ZN => n9136);
   U14669 : OAI22_X1 port map( A1 => n1436_port, A2 => n10636, B1 => n1372_port
                           , B2 => n10627, ZN => n9154);
   U14670 : OAI22_X1 port map( A1 => n1435_port, A2 => n10636, B1 => n1371_port
                           , B2 => n10627, ZN => n9172);
   U14671 : OAI22_X1 port map( A1 => n1434_port, A2 => n10636, B1 => n1370_port
                           , B2 => n10627, ZN => n9190);
   U14672 : OAI22_X1 port map( A1 => n1433_port, A2 => n10636, B1 => n1369_port
                           , B2 => n10627, ZN => n9208);
   U14673 : OAI22_X1 port map( A1 => n1432_port, A2 => n10635, B1 => n1368_port
                           , B2 => n10626, ZN => n9226);
   U14674 : OAI22_X1 port map( A1 => n1431_port, A2 => n10635, B1 => n1367_port
                           , B2 => n10626, ZN => n9244);
   U14675 : OAI22_X1 port map( A1 => n1430_port, A2 => n10635, B1 => n1366_port
                           , B2 => n10626, ZN => n9262);
   U14676 : OAI22_X1 port map( A1 => n1429_port, A2 => n10635, B1 => n1365_port
                           , B2 => n10626, ZN => n9280);
   U14677 : OAI22_X1 port map( A1 => n1428_port, A2 => n10635, B1 => n1364_port
                           , B2 => n10626, ZN => n9298);
   U14678 : OAI22_X1 port map( A1 => n1427_port, A2 => n10635, B1 => n1363_port
                           , B2 => n10626, ZN => n9316);
   U14679 : OAI22_X1 port map( A1 => n1426_port, A2 => n10635, B1 => n1362_port
                           , B2 => n10626, ZN => n9334);
   U14680 : OAI22_X1 port map( A1 => n1425_port, A2 => n10635, B1 => n1361_port
                           , B2 => n10626, ZN => n9352);
   U14681 : OAI22_X1 port map( A1 => n1424_port, A2 => n10635, B1 => n1360_port
                           , B2 => n10626, ZN => n9370);
   U14682 : OAI22_X1 port map( A1 => n1423_port, A2 => n10635, B1 => n1359_port
                           , B2 => n10626, ZN => n9388);
   U14683 : OAI22_X1 port map( A1 => n1422_port, A2 => n10635, B1 => n1358_port
                           , B2 => n10626, ZN => n9406);
   U14684 : OAI22_X1 port map( A1 => n1421_port, A2 => n10635, B1 => n1357_port
                           , B2 => n10626, ZN => n9424);
   U14685 : OAI22_X1 port map( A1 => n1420_port, A2 => n10634, B1 => n1356_port
                           , B2 => n10625, ZN => n9442);
   U14686 : OAI22_X1 port map( A1 => n1419_port, A2 => n10634, B1 => n1355_port
                           , B2 => n10625, ZN => n9460);
   U14687 : OAI22_X1 port map( A1 => n1418_port, A2 => n10634, B1 => n1354_port
                           , B2 => n10625, ZN => n9478);
   U14688 : OAI22_X1 port map( A1 => n1417_port, A2 => n10634, B1 => n1353_port
                           , B2 => n10625, ZN => n9496);
   U14689 : OAI22_X1 port map( A1 => n1416_port, A2 => n10634, B1 => n1352_port
                           , B2 => n10625, ZN => n9514);
   U14690 : OAI22_X1 port map( A1 => n1415_port, A2 => n10634, B1 => n1351_port
                           , B2 => n10625, ZN => n9532);
   U14691 : OAI22_X1 port map( A1 => n1414_port, A2 => n10634, B1 => n1350_port
                           , B2 => n10625, ZN => n9550);
   U14692 : OAI22_X1 port map( A1 => n1413_port, A2 => n10634, B1 => n1349_port
                           , B2 => n10625, ZN => n9568);
   U14693 : OAI22_X1 port map( A1 => n1412_port, A2 => n10634, B1 => n1348_port
                           , B2 => n10625, ZN => n9586);
   U14694 : OAI22_X1 port map( A1 => n1411_port, A2 => n10634, B1 => n1347_port
                           , B2 => n10625, ZN => n9604);
   U14695 : OAI22_X1 port map( A1 => n1410_port, A2 => n10634, B1 => n1346_port
                           , B2 => n10625, ZN => n9622);
   U14696 : OAI22_X1 port map( A1 => n1409_port, A2 => n10634, B1 => n1345_port
                           , B2 => n10625, ZN => n9646);
   U14697 : OAI22_X1 port map( A1 => n2048_port, A2 => n10983, B1 => n1984_port
                           , B2 => n10974, ZN => n7291);
   U14698 : OAI22_X1 port map( A1 => n2047_port, A2 => n10983, B1 => n1983_port
                           , B2 => n10974, ZN => n7331);
   U14699 : OAI22_X1 port map( A1 => n2046_port, A2 => n10983, B1 => n1982_port
                           , B2 => n10974, ZN => n7349);
   U14700 : OAI22_X1 port map( A1 => n2045_port, A2 => n10983, B1 => n1981_port
                           , B2 => n10974, ZN => n7367);
   U14701 : OAI22_X1 port map( A1 => n2044_port, A2 => n10982, B1 => n1980_port
                           , B2 => n10973, ZN => n7385);
   U14702 : OAI22_X1 port map( A1 => n2043_port, A2 => n10982, B1 => n1979_port
                           , B2 => n10973, ZN => n7403);
   U14703 : OAI22_X1 port map( A1 => n2042_port, A2 => n10982, B1 => n1978_port
                           , B2 => n10973, ZN => n7421);
   U14704 : OAI22_X1 port map( A1 => n2041_port, A2 => n10982, B1 => n1977_port
                           , B2 => n10973, ZN => n7439);
   U14705 : OAI22_X1 port map( A1 => n2040_port, A2 => n10982, B1 => n1976_port
                           , B2 => n10973, ZN => n7457);
   U14706 : OAI22_X1 port map( A1 => n2039_port, A2 => n10982, B1 => n1975_port
                           , B2 => n10973, ZN => n7475);
   U14707 : OAI22_X1 port map( A1 => n2038_port, A2 => n10982, B1 => n1974_port
                           , B2 => n10973, ZN => n7493);
   U14708 : OAI22_X1 port map( A1 => n2037_port, A2 => n10982, B1 => n1973_port
                           , B2 => n10973, ZN => n7511);
   U14709 : OAI22_X1 port map( A1 => n2036_port, A2 => n10982, B1 => n1972_port
                           , B2 => n10973, ZN => n7529);
   U14710 : OAI22_X1 port map( A1 => n2035_port, A2 => n10982, B1 => n1971_port
                           , B2 => n10973, ZN => n7547);
   U14711 : OAI22_X1 port map( A1 => n2034_port, A2 => n10982, B1 => n1970_port
                           , B2 => n10973, ZN => n7565);
   U14712 : OAI22_X1 port map( A1 => n2033_port, A2 => n10982, B1 => n1969_port
                           , B2 => n10973, ZN => n7583);
   U14713 : OAI22_X1 port map( A1 => n2032_port, A2 => n10981, B1 => n1968_port
                           , B2 => n10972, ZN => n7601);
   U14714 : OAI22_X1 port map( A1 => n2031_port, A2 => n10981, B1 => n1967_port
                           , B2 => n10972, ZN => n7619);
   U14715 : OAI22_X1 port map( A1 => n2030_port, A2 => n10981, B1 => n1966_port
                           , B2 => n10972, ZN => n7637);
   U14716 : OAI22_X1 port map( A1 => n2029_port, A2 => n10981, B1 => n1965_port
                           , B2 => n10972, ZN => n7655);
   U14717 : OAI22_X1 port map( A1 => n2028_port, A2 => n10981, B1 => n1964_port
                           , B2 => n10972, ZN => n7673);
   U14718 : OAI22_X1 port map( A1 => n2027_port, A2 => n10981, B1 => n1963_port
                           , B2 => n10972, ZN => n7691);
   U14719 : OAI22_X1 port map( A1 => n2026_port, A2 => n10981, B1 => n1962_port
                           , B2 => n10972, ZN => n7709);
   U14720 : OAI22_X1 port map( A1 => n2025_port, A2 => n10981, B1 => n1961_port
                           , B2 => n10972, ZN => n7727);
   U14721 : OAI22_X1 port map( A1 => n2024_port, A2 => n10981, B1 => n1960_port
                           , B2 => n10972, ZN => n7745);
   U14722 : OAI22_X1 port map( A1 => n2023_port, A2 => n10981, B1 => n1959_port
                           , B2 => n10972, ZN => n7763);
   U14723 : OAI22_X1 port map( A1 => n2022_port, A2 => n10981, B1 => n1958_port
                           , B2 => n10972, ZN => n7781);
   U14724 : OAI22_X1 port map( A1 => n2021_port, A2 => n10981, B1 => n1957_port
                           , B2 => n10972, ZN => n7799);
   U14725 : OAI22_X1 port map( A1 => n2020_port, A2 => n10980, B1 => n1956_port
                           , B2 => n10971, ZN => n7817);
   U14726 : OAI22_X1 port map( A1 => n2019_port, A2 => n10980, B1 => n1955_port
                           , B2 => n10971, ZN => n7835);
   U14727 : OAI22_X1 port map( A1 => n2018_port, A2 => n10980, B1 => n1954_port
                           , B2 => n10971, ZN => n7853);
   U14728 : OAI22_X1 port map( A1 => n2017_port, A2 => n10980, B1 => n1953_port
                           , B2 => n10971, ZN => n7871);
   U14729 : OAI22_X1 port map( A1 => n2016_port, A2 => n10980, B1 => n1952_port
                           , B2 => n10971, ZN => n7889);
   U14730 : OAI22_X1 port map( A1 => n2015_port, A2 => n10980, B1 => n1951_port
                           , B2 => n10971, ZN => n7907);
   U14731 : OAI22_X1 port map( A1 => n2014_port, A2 => n10980, B1 => n1950_port
                           , B2 => n10971, ZN => n7925);
   U14732 : OAI22_X1 port map( A1 => n2013_port, A2 => n10980, B1 => n1949_port
                           , B2 => n10971, ZN => n7943);
   U14733 : OAI22_X1 port map( A1 => n2012_port, A2 => n10980, B1 => n1948_port
                           , B2 => n10971, ZN => n7961);
   U14734 : OAI22_X1 port map( A1 => n2011_port, A2 => n10980, B1 => n1947_port
                           , B2 => n10971, ZN => n7979);
   U14735 : OAI22_X1 port map( A1 => n2010_port, A2 => n10980, B1 => n1946_port
                           , B2 => n10971, ZN => n7997);
   U14736 : OAI22_X1 port map( A1 => n2009_port, A2 => n10980, B1 => n1945_port
                           , B2 => n10971, ZN => n8015);
   U14737 : OAI22_X1 port map( A1 => n2008_port, A2 => n10979, B1 => n1944_port
                           , B2 => n10970, ZN => n8033);
   U14738 : OAI22_X1 port map( A1 => n2007_port, A2 => n10979, B1 => n1943_port
                           , B2 => n10970, ZN => n8051);
   U14739 : OAI22_X1 port map( A1 => n2006_port, A2 => n10979, B1 => n1942_port
                           , B2 => n10970, ZN => n8069);
   U14740 : OAI22_X1 port map( A1 => n2005_port, A2 => n10979, B1 => n1941_port
                           , B2 => n10970, ZN => n8087);
   U14741 : OAI22_X1 port map( A1 => n2004_port, A2 => n10979, B1 => n1940_port
                           , B2 => n10970, ZN => n8105);
   U14742 : OAI22_X1 port map( A1 => n2003_port, A2 => n10979, B1 => n1939_port
                           , B2 => n10970, ZN => n8123);
   U14743 : OAI22_X1 port map( A1 => n2002_port, A2 => n10979, B1 => n1938_port
                           , B2 => n10970, ZN => n8141);
   U14744 : OAI22_X1 port map( A1 => n2001_port, A2 => n10979, B1 => n1937_port
                           , B2 => n10970, ZN => n8159);
   U14745 : OAI22_X1 port map( A1 => n2000_port, A2 => n10979, B1 => n1936_port
                           , B2 => n10970, ZN => n8177);
   U14746 : OAI22_X1 port map( A1 => n1999_port, A2 => n10979, B1 => n1935_port
                           , B2 => n10970, ZN => n8195);
   U14747 : OAI22_X1 port map( A1 => n1998_port, A2 => n10979, B1 => n1934_port
                           , B2 => n10970, ZN => n8213);
   U14748 : OAI22_X1 port map( A1 => n1997_port, A2 => n10979, B1 => n1933_port
                           , B2 => n10970, ZN => n8231);
   U14749 : OAI22_X1 port map( A1 => n1996_port, A2 => n10978, B1 => n1932_port
                           , B2 => n10969, ZN => n8249);
   U14750 : OAI22_X1 port map( A1 => n1995_port, A2 => n10978, B1 => n1931_port
                           , B2 => n10969, ZN => n8267);
   U14751 : OAI22_X1 port map( A1 => n1994_port, A2 => n10978, B1 => n1930_port
                           , B2 => n10969, ZN => n8285);
   U14752 : OAI22_X1 port map( A1 => n1993_port, A2 => n10978, B1 => n1929_port
                           , B2 => n10969, ZN => n8303);
   U14753 : OAI22_X1 port map( A1 => n1992_port, A2 => n10978, B1 => n1928_port
                           , B2 => n10969, ZN => n8321);
   U14754 : OAI22_X1 port map( A1 => n1991_port, A2 => n10978, B1 => n1927_port
                           , B2 => n10969, ZN => n8339);
   U14755 : OAI22_X1 port map( A1 => n1990_port, A2 => n10978, B1 => n1926_port
                           , B2 => n10969, ZN => n8357);
   U14756 : OAI22_X1 port map( A1 => n1989_port, A2 => n10978, B1 => n1925_port
                           , B2 => n10969, ZN => n8375);
   U14757 : OAI22_X1 port map( A1 => n1988_port, A2 => n10978, B1 => n1924_port
                           , B2 => n10969, ZN => n8393);
   U14758 : OAI22_X1 port map( A1 => n1987_port, A2 => n10978, B1 => n1923_port
                           , B2 => n10969, ZN => n8411);
   U14759 : OAI22_X1 port map( A1 => n1986_port, A2 => n10978, B1 => n1922_port
                           , B2 => n10969, ZN => n8429);
   U14760 : OAI22_X1 port map( A1 => n1985_port, A2 => n10978, B1 => n1921_port
                           , B2 => n10969, ZN => n8447);
   U14761 : OAI22_X1 port map( A1 => n2048_port, A2 => n10758, B1 => n1984_port
                           , B2 => n10749, ZN => n8471);
   U14762 : OAI22_X1 port map( A1 => n2047_port, A2 => n10758, B1 => n1983_port
                           , B2 => n10749, ZN => n8511);
   U14763 : OAI22_X1 port map( A1 => n2046_port, A2 => n10758, B1 => n1982_port
                           , B2 => n10749, ZN => n8529);
   U14764 : OAI22_X1 port map( A1 => n2045_port, A2 => n10758, B1 => n1981_port
                           , B2 => n10749, ZN => n8547);
   U14765 : OAI22_X1 port map( A1 => n2044_port, A2 => n10757, B1 => n1980_port
                           , B2 => n10748, ZN => n8565);
   U14766 : OAI22_X1 port map( A1 => n2043_port, A2 => n10757, B1 => n1979_port
                           , B2 => n10748, ZN => n8583);
   U14767 : OAI22_X1 port map( A1 => n2042_port, A2 => n10757, B1 => n1978_port
                           , B2 => n10748, ZN => n8601);
   U14768 : OAI22_X1 port map( A1 => n2041_port, A2 => n10757, B1 => n1977_port
                           , B2 => n10748, ZN => n8619);
   U14769 : OAI22_X1 port map( A1 => n2040_port, A2 => n10757, B1 => n1976_port
                           , B2 => n10748, ZN => n8637);
   U14770 : OAI22_X1 port map( A1 => n2039_port, A2 => n10757, B1 => n1975_port
                           , B2 => n10748, ZN => n8655);
   U14771 : OAI22_X1 port map( A1 => n2038_port, A2 => n10757, B1 => n1974_port
                           , B2 => n10748, ZN => n8673);
   U14772 : OAI22_X1 port map( A1 => n2037_port, A2 => n10757, B1 => n1973_port
                           , B2 => n10748, ZN => n8691);
   U14773 : OAI22_X1 port map( A1 => n2036_port, A2 => n10757, B1 => n1972_port
                           , B2 => n10748, ZN => n8709);
   U14774 : OAI22_X1 port map( A1 => n2035_port, A2 => n10757, B1 => n1971_port
                           , B2 => n10748, ZN => n8727);
   U14775 : OAI22_X1 port map( A1 => n2034_port, A2 => n10757, B1 => n1970_port
                           , B2 => n10748, ZN => n8745);
   U14776 : OAI22_X1 port map( A1 => n2033_port, A2 => n10757, B1 => n1969_port
                           , B2 => n10748, ZN => n8763);
   U14777 : OAI22_X1 port map( A1 => n2032_port, A2 => n10756, B1 => n1968_port
                           , B2 => n10747, ZN => n8781);
   U14778 : OAI22_X1 port map( A1 => n2031_port, A2 => n10756, B1 => n1967_port
                           , B2 => n10747, ZN => n8799);
   U14779 : OAI22_X1 port map( A1 => n2030_port, A2 => n10756, B1 => n1966_port
                           , B2 => n10747, ZN => n8817);
   U14780 : OAI22_X1 port map( A1 => n2029_port, A2 => n10756, B1 => n1965_port
                           , B2 => n10747, ZN => n8835);
   U14781 : OAI22_X1 port map( A1 => n2028_port, A2 => n10756, B1 => n1964_port
                           , B2 => n10747, ZN => n8853);
   U14782 : OAI22_X1 port map( A1 => n2027_port, A2 => n10756, B1 => n1963_port
                           , B2 => n10747, ZN => n8871);
   U14783 : OAI22_X1 port map( A1 => n2026_port, A2 => n10756, B1 => n1962_port
                           , B2 => n10747, ZN => n8889);
   U14784 : OAI22_X1 port map( A1 => n2025_port, A2 => n10756, B1 => n1961_port
                           , B2 => n10747, ZN => n8907);
   U14785 : OAI22_X1 port map( A1 => n2024_port, A2 => n10756, B1 => n1960_port
                           , B2 => n10747, ZN => n8925);
   U14786 : OAI22_X1 port map( A1 => n2023_port, A2 => n10756, B1 => n1959_port
                           , B2 => n10747, ZN => n8943);
   U14787 : OAI22_X1 port map( A1 => n2022_port, A2 => n10756, B1 => n1958_port
                           , B2 => n10747, ZN => n8961);
   U14788 : OAI22_X1 port map( A1 => n2021_port, A2 => n10756, B1 => n1957_port
                           , B2 => n10747, ZN => n8979);
   U14789 : OAI22_X1 port map( A1 => n2020_port, A2 => n10755, B1 => n1956_port
                           , B2 => n10746, ZN => n8997);
   U14790 : OAI22_X1 port map( A1 => n2019_port, A2 => n10755, B1 => n1955_port
                           , B2 => n10746, ZN => n9015);
   U14791 : OAI22_X1 port map( A1 => n2018_port, A2 => n10755, B1 => n1954_port
                           , B2 => n10746, ZN => n9033);
   U14792 : OAI22_X1 port map( A1 => n2017_port, A2 => n10755, B1 => n1953_port
                           , B2 => n10746, ZN => n9051);
   U14793 : OAI22_X1 port map( A1 => n2016_port, A2 => n10755, B1 => n1952_port
                           , B2 => n10746, ZN => n9069);
   U14794 : OAI22_X1 port map( A1 => n2015_port, A2 => n10755, B1 => n1951_port
                           , B2 => n10746, ZN => n9087);
   U14795 : OAI22_X1 port map( A1 => n2014_port, A2 => n10755, B1 => n1950_port
                           , B2 => n10746, ZN => n9105);
   U14796 : OAI22_X1 port map( A1 => n2013_port, A2 => n10755, B1 => n1949_port
                           , B2 => n10746, ZN => n9123);
   U14797 : OAI22_X1 port map( A1 => n2012_port, A2 => n10755, B1 => n1948_port
                           , B2 => n10746, ZN => n9141);
   U14798 : OAI22_X1 port map( A1 => n2011_port, A2 => n10755, B1 => n1947_port
                           , B2 => n10746, ZN => n9159);
   U14799 : OAI22_X1 port map( A1 => n2010_port, A2 => n10755, B1 => n1946_port
                           , B2 => n10746, ZN => n9177);
   U14800 : OAI22_X1 port map( A1 => n2009_port, A2 => n10755, B1 => n1945_port
                           , B2 => n10746, ZN => n9195);
   U14801 : OAI22_X1 port map( A1 => n2008_port, A2 => n10754, B1 => n1944_port
                           , B2 => n10745, ZN => n9213);
   U14802 : OAI22_X1 port map( A1 => n2007_port, A2 => n10754, B1 => n1943_port
                           , B2 => n10745, ZN => n9231);
   U14803 : OAI22_X1 port map( A1 => n2006_port, A2 => n10754, B1 => n1942_port
                           , B2 => n10745, ZN => n9249);
   U14804 : OAI22_X1 port map( A1 => n2005_port, A2 => n10754, B1 => n1941_port
                           , B2 => n10745, ZN => n9267);
   U14805 : OAI22_X1 port map( A1 => n2004_port, A2 => n10754, B1 => n1940_port
                           , B2 => n10745, ZN => n9285);
   U14806 : OAI22_X1 port map( A1 => n2003_port, A2 => n10754, B1 => n1939_port
                           , B2 => n10745, ZN => n9303);
   U14807 : OAI22_X1 port map( A1 => n2002_port, A2 => n10754, B1 => n1938_port
                           , B2 => n10745, ZN => n9321);
   U14808 : OAI22_X1 port map( A1 => n2001_port, A2 => n10754, B1 => n1937_port
                           , B2 => n10745, ZN => n9339);
   U14809 : OAI22_X1 port map( A1 => n2000_port, A2 => n10754, B1 => n1936_port
                           , B2 => n10745, ZN => n9357);
   U14810 : OAI22_X1 port map( A1 => n1999_port, A2 => n10754, B1 => n1935_port
                           , B2 => n10745, ZN => n9375);
   U14811 : OAI22_X1 port map( A1 => n1998_port, A2 => n10754, B1 => n1934_port
                           , B2 => n10745, ZN => n9393);
   U14812 : OAI22_X1 port map( A1 => n1997_port, A2 => n10754, B1 => n1933_port
                           , B2 => n10745, ZN => n9411);
   U14813 : OAI22_X1 port map( A1 => n1996_port, A2 => n10753, B1 => n1932_port
                           , B2 => n10744, ZN => n9429);
   U14814 : OAI22_X1 port map( A1 => n1995_port, A2 => n10753, B1 => n1931_port
                           , B2 => n10744, ZN => n9447);
   U14815 : OAI22_X1 port map( A1 => n1994_port, A2 => n10753, B1 => n1930_port
                           , B2 => n10744, ZN => n9465);
   U14816 : OAI22_X1 port map( A1 => n1993_port, A2 => n10753, B1 => n1929_port
                           , B2 => n10744, ZN => n9483);
   U14817 : OAI22_X1 port map( A1 => n1992_port, A2 => n10753, B1 => n1928_port
                           , B2 => n10744, ZN => n9501);
   U14818 : OAI22_X1 port map( A1 => n1991_port, A2 => n10753, B1 => n1927_port
                           , B2 => n10744, ZN => n9519);
   U14819 : OAI22_X1 port map( A1 => n1990_port, A2 => n10753, B1 => n1926_port
                           , B2 => n10744, ZN => n9537);
   U14820 : OAI22_X1 port map( A1 => n1989_port, A2 => n10753, B1 => n1925_port
                           , B2 => n10744, ZN => n9555);
   U14821 : OAI22_X1 port map( A1 => n1988_port, A2 => n10753, B1 => n1924_port
                           , B2 => n10744, ZN => n9573);
   U14822 : OAI22_X1 port map( A1 => n1987_port, A2 => n10753, B1 => n1923_port
                           , B2 => n10744, ZN => n9591);
   U14823 : OAI22_X1 port map( A1 => n1986_port, A2 => n10753, B1 => n1922_port
                           , B2 => n10744, ZN => n9609);
   U14824 : OAI22_X1 port map( A1 => n1985_port, A2 => n10753, B1 => n1921_port
                           , B2 => n10744, ZN => n9627);
   U14825 : AOI21_X1 port map( B1 => n7294, B2 => n7295, A => n11071, ZN => 
                           n7293);
   U14826 : AOI221_X1 port map( B1 => n11017, B2 => n10287, C1 => n11000, C2 =>
                           n9839, A => n7302, ZN => n7294);
   U14827 : AOI221_X1 port map( B1 => n11052, B2 => n10288, C1 => n11029, C2 =>
                           n9840, A => n7299, ZN => n7295);
   U14828 : OAI22_X1 port map( A1 => n128_port, A2 => n11594, B1 => n256_port, 
                           B2 => n11577, ZN => n7302);
   U14829 : AOI21_X1 port map( B1 => n7334, B2 => n7335, A => n11071, ZN => 
                           n7333);
   U14830 : AOI221_X1 port map( B1 => n11012, B2 => n10289, C1 => n10995, C2 =>
                           n9841, A => n7337, ZN => n7334);
   U14831 : AOI221_X1 port map( B1 => n11047, B2 => n10290, C1 => n11029, C2 =>
                           n9842, A => n7336, ZN => n7335);
   U14832 : OAI22_X1 port map( A1 => n127_port, A2 => n11594, B1 => n255_port, 
                           B2 => n11577, ZN => n7337);
   U14833 : AOI21_X1 port map( B1 => n7352, B2 => n7353, A => n11071, ZN => 
                           n7351);
   U14834 : AOI221_X1 port map( B1 => n11012, B2 => n10291, C1 => n10995, C2 =>
                           n9843, A => n7355, ZN => n7352);
   U14835 : AOI221_X1 port map( B1 => n11047, B2 => n10292, C1 => n11029, C2 =>
                           n9844, A => n7354, ZN => n7353);
   U14836 : OAI22_X1 port map( A1 => n126_port, A2 => n11594, B1 => n254_port, 
                           B2 => n11577, ZN => n7355);
   U14837 : AOI21_X1 port map( B1 => n7370, B2 => n7371, A => n11071, ZN => 
                           n7369);
   U14838 : AOI221_X1 port map( B1 => n11012, B2 => n10293, C1 => n10995, C2 =>
                           n9845, A => n7373, ZN => n7370);
   U14839 : AOI221_X1 port map( B1 => n11047, B2 => n10294, C1 => n11029, C2 =>
                           n9846, A => n7372, ZN => n7371);
   U14840 : OAI22_X1 port map( A1 => n125_port, A2 => n11594, B1 => n253_port, 
                           B2 => n11577, ZN => n7373);
   U14841 : AOI21_X1 port map( B1 => n7388, B2 => n7389, A => n11070, ZN => 
                           n7387);
   U14842 : AOI221_X1 port map( B1 => n11012, B2 => n10295, C1 => n10995, C2 =>
                           n9847, A => n7391, ZN => n7388);
   U14843 : AOI221_X1 port map( B1 => n11047, B2 => n10296, C1 => n11029, C2 =>
                           n9848, A => n7390, ZN => n7389);
   U14844 : OAI22_X1 port map( A1 => n124_port, A2 => n11593, B1 => n252_port, 
                           B2 => n11576, ZN => n7391);
   U14845 : AOI21_X1 port map( B1 => n7406, B2 => n7407, A => n11070, ZN => 
                           n7405);
   U14846 : AOI221_X1 port map( B1 => n11012, B2 => n10297, C1 => n10995, C2 =>
                           n9849, A => n7409, ZN => n7406);
   U14847 : AOI221_X1 port map( B1 => n11047, B2 => n10298, C1 => n11029, C2 =>
                           n9850, A => n7408, ZN => n7407);
   U14848 : OAI22_X1 port map( A1 => n123_port, A2 => n11593, B1 => n251_port, 
                           B2 => n11576, ZN => n7409);
   U14849 : AOI21_X1 port map( B1 => n7424, B2 => n7425, A => n11070, ZN => 
                           n7423);
   U14850 : AOI221_X1 port map( B1 => n11012, B2 => n10299, C1 => n10995, C2 =>
                           n9851, A => n7427, ZN => n7424);
   U14851 : AOI221_X1 port map( B1 => n11047, B2 => n10300, C1 => n11030, C2 =>
                           n9852, A => n7426, ZN => n7425);
   U14852 : OAI22_X1 port map( A1 => n122_port, A2 => n11593, B1 => n250_port, 
                           B2 => n11576, ZN => n7427);
   U14853 : AOI21_X1 port map( B1 => n7442, B2 => n7443, A => n11070, ZN => 
                           n7441);
   U14854 : AOI221_X1 port map( B1 => n11013, B2 => n10301, C1 => n10996, C2 =>
                           n9853, A => n7445, ZN => n7442);
   U14855 : AOI221_X1 port map( B1 => n11048, B2 => n10302, C1 => n11030, C2 =>
                           n9854, A => n7444, ZN => n7443);
   U14856 : OAI22_X1 port map( A1 => n121_port, A2 => n11593, B1 => n249_port, 
                           B2 => n11576, ZN => n7445);
   U14857 : AOI21_X1 port map( B1 => n7460, B2 => n7461, A => n11070, ZN => 
                           n7459);
   U14858 : AOI221_X1 port map( B1 => n11013, B2 => n10303, C1 => n10996, C2 =>
                           n9855, A => n7463, ZN => n7460);
   U14859 : AOI221_X1 port map( B1 => n11048, B2 => n10304, C1 => n11030, C2 =>
                           n9856, A => n7462, ZN => n7461);
   U14860 : OAI22_X1 port map( A1 => n120_port, A2 => n11593, B1 => n248_port, 
                           B2 => n11576, ZN => n7463);
   U14861 : AOI21_X1 port map( B1 => n7478, B2 => n7479, A => n11070, ZN => 
                           n7477);
   U14862 : AOI221_X1 port map( B1 => n11013, B2 => n10305, C1 => n10996, C2 =>
                           n9857, A => n7481, ZN => n7478);
   U14863 : AOI221_X1 port map( B1 => n11048, B2 => n10306, C1 => n11030, C2 =>
                           n9858, A => n7480, ZN => n7479);
   U14864 : OAI22_X1 port map( A1 => n119_port, A2 => n11593, B1 => n247_port, 
                           B2 => n11576, ZN => n7481);
   U14865 : AOI21_X1 port map( B1 => n7496, B2 => n7497, A => n11070, ZN => 
                           n7495);
   U14866 : AOI221_X1 port map( B1 => n11013, B2 => n10307, C1 => n10996, C2 =>
                           n9859, A => n7499, ZN => n7496);
   U14867 : AOI221_X1 port map( B1 => n11048, B2 => n10308, C1 => n11030, C2 =>
                           n9860, A => n7498, ZN => n7497);
   U14868 : OAI22_X1 port map( A1 => n118_port, A2 => n11592, B1 => n246_port, 
                           B2 => n11575, ZN => n7499);
   U14869 : AOI21_X1 port map( B1 => n7514, B2 => n7515, A => n11070, ZN => 
                           n7513);
   U14870 : AOI221_X1 port map( B1 => n11013, B2 => n10309, C1 => n10996, C2 =>
                           n9861, A => n7517, ZN => n7514);
   U14871 : AOI221_X1 port map( B1 => n11048, B2 => n10310, C1 => n11030, C2 =>
                           n9862, A => n7516, ZN => n7515);
   U14872 : OAI22_X1 port map( A1 => n117_port, A2 => n11592, B1 => n245_port, 
                           B2 => n11575, ZN => n7517);
   U14873 : AOI21_X1 port map( B1 => n7532, B2 => n7533, A => n11070, ZN => 
                           n7531);
   U14874 : AOI221_X1 port map( B1 => n11013, B2 => n10311, C1 => n10996, C2 =>
                           n9863, A => n7535, ZN => n7532);
   U14875 : AOI221_X1 port map( B1 => n11048, B2 => n10312, C1 => n11031, C2 =>
                           n9864, A => n7534, ZN => n7533);
   U14876 : OAI22_X1 port map( A1 => n116_port, A2 => n11592, B1 => n244_port, 
                           B2 => n11575, ZN => n7535);
   U14877 : AOI21_X1 port map( B1 => n7550, B2 => n7551, A => n11070, ZN => 
                           n7549);
   U14878 : AOI221_X1 port map( B1 => n11014, B2 => n10313, C1 => n10997, C2 =>
                           n9865, A => n7553, ZN => n7550);
   U14879 : AOI221_X1 port map( B1 => n11049, B2 => n10314, C1 => n11031, C2 =>
                           n9866, A => n7552, ZN => n7551);
   U14880 : OAI22_X1 port map( A1 => n115_port, A2 => n11592, B1 => n243_port, 
                           B2 => n11575, ZN => n7553);
   U14881 : AOI21_X1 port map( B1 => n7568, B2 => n7569, A => n11070, ZN => 
                           n7567);
   U14882 : AOI221_X1 port map( B1 => n11014, B2 => n10315, C1 => n10997, C2 =>
                           n9867, A => n7571, ZN => n7568);
   U14883 : AOI221_X1 port map( B1 => n11049, B2 => n10316, C1 => n11031, C2 =>
                           n9868, A => n7570, ZN => n7569);
   U14884 : OAI22_X1 port map( A1 => n114_port, A2 => n11592, B1 => n242_port, 
                           B2 => n11575, ZN => n7571);
   U14885 : AOI21_X1 port map( B1 => n7586, B2 => n7587, A => n11070, ZN => 
                           n7585);
   U14886 : AOI221_X1 port map( B1 => n11014, B2 => n10317, C1 => n10997, C2 =>
                           n9869, A => n7589, ZN => n7586);
   U14887 : AOI221_X1 port map( B1 => n11049, B2 => n10318, C1 => n11031, C2 =>
                           n9870, A => n7588, ZN => n7587);
   U14888 : OAI22_X1 port map( A1 => n113_port, A2 => n11592, B1 => n241_port, 
                           B2 => n11575, ZN => n7589);
   U14889 : AOI21_X1 port map( B1 => n7604, B2 => n7605, A => n11069, ZN => 
                           n7603);
   U14890 : AOI221_X1 port map( B1 => n11014, B2 => n10319, C1 => n10997, C2 =>
                           n9871, A => n7607, ZN => n7604);
   U14891 : AOI221_X1 port map( B1 => n11049, B2 => n10320, C1 => n11031, C2 =>
                           n9872, A => n7606, ZN => n7605);
   U14892 : OAI22_X1 port map( A1 => n112_port, A2 => n11591, B1 => n240_port, 
                           B2 => n11574, ZN => n7607);
   U14893 : AOI21_X1 port map( B1 => n7622, B2 => n7623, A => n11069, ZN => 
                           n7621);
   U14894 : AOI221_X1 port map( B1 => n11014, B2 => n10321, C1 => n10997, C2 =>
                           n9873, A => n7625, ZN => n7622);
   U14895 : AOI221_X1 port map( B1 => n11049, B2 => n10322, C1 => n11031, C2 =>
                           n9874, A => n7624, ZN => n7623);
   U14896 : OAI22_X1 port map( A1 => n111_port, A2 => n11591, B1 => n239_port, 
                           B2 => n11574, ZN => n7625);
   U14897 : AOI21_X1 port map( B1 => n7640, B2 => n7641, A => n11069, ZN => 
                           n7639);
   U14898 : AOI221_X1 port map( B1 => n11014, B2 => n10323, C1 => n10997, C2 =>
                           n9875, A => n7643, ZN => n7640);
   U14899 : AOI221_X1 port map( B1 => n11049, B2 => n10324, C1 => n11032, C2 =>
                           n9876, A => n7642, ZN => n7641);
   U14900 : OAI22_X1 port map( A1 => n110_port, A2 => n11591, B1 => n238_port, 
                           B2 => n11574, ZN => n7643);
   U14901 : AOI21_X1 port map( B1 => n7658, B2 => n7659, A => n11069, ZN => 
                           n7657);
   U14902 : AOI221_X1 port map( B1 => n11014, B2 => n10325, C1 => n10997, C2 =>
                           n9877, A => n7661, ZN => n7658);
   U14903 : AOI221_X1 port map( B1 => n11050, B2 => n10326, C1 => n11032, C2 =>
                           n9878, A => n7660, ZN => n7659);
   U14904 : OAI22_X1 port map( A1 => n109_port, A2 => n11591, B1 => n237_port, 
                           B2 => n11574, ZN => n7661);
   U14905 : AOI21_X1 port map( B1 => n7676, B2 => n7677, A => n11069, ZN => 
                           n7675);
   U14906 : AOI221_X1 port map( B1 => n11015, B2 => n10327, C1 => n10998, C2 =>
                           n9879, A => n7679, ZN => n7676);
   U14907 : AOI221_X1 port map( B1 => n11050, B2 => n10328, C1 => n11032, C2 =>
                           n9880, A => n7678, ZN => n7677);
   U14908 : OAI22_X1 port map( A1 => n108_port, A2 => n11591, B1 => n236_port, 
                           B2 => n11574, ZN => n7679);
   U14909 : AOI21_X1 port map( B1 => n7694, B2 => n7695, A => n11069, ZN => 
                           n7693);
   U14910 : AOI221_X1 port map( B1 => n11015, B2 => n10329, C1 => n10998, C2 =>
                           n9881, A => n7697, ZN => n7694);
   U14911 : AOI221_X1 port map( B1 => n11050, B2 => n10330, C1 => n11032, C2 =>
                           n9882, A => n7696, ZN => n7695);
   U14912 : OAI22_X1 port map( A1 => n107_port, A2 => n11591, B1 => n235_port, 
                           B2 => n11574, ZN => n7697);
   U14913 : AOI21_X1 port map( B1 => n7712, B2 => n7713, A => n11069, ZN => 
                           n7711);
   U14914 : AOI221_X1 port map( B1 => n11015, B2 => n10331, C1 => n10998, C2 =>
                           n9883, A => n7715, ZN => n7712);
   U14915 : AOI221_X1 port map( B1 => n11050, B2 => n10332, C1 => n11032, C2 =>
                           n9884, A => n7714, ZN => n7713);
   U14916 : OAI22_X1 port map( A1 => n106_port, A2 => n11590, B1 => n234_port, 
                           B2 => n11573, ZN => n7715);
   U14917 : AOI21_X1 port map( B1 => n7730, B2 => n7731, A => n11069, ZN => 
                           n7729);
   U14918 : AOI221_X1 port map( B1 => n11015, B2 => n10333, C1 => n10998, C2 =>
                           n9885, A => n7733, ZN => n7730);
   U14919 : AOI221_X1 port map( B1 => n11050, B2 => n10334, C1 => n11032, C2 =>
                           n9886, A => n7732, ZN => n7731);
   U14920 : OAI22_X1 port map( A1 => n105_port, A2 => n11590, B1 => n233_port, 
                           B2 => n11573, ZN => n7733);
   U14921 : AOI21_X1 port map( B1 => n7748, B2 => n7749, A => n11069, ZN => 
                           n7747);
   U14922 : AOI221_X1 port map( B1 => n11015, B2 => n10335, C1 => n10998, C2 =>
                           n9887, A => n7751, ZN => n7748);
   U14923 : AOI221_X1 port map( B1 => n11050, B2 => n10336, C1 => n11033, C2 =>
                           n9888, A => n7750, ZN => n7749);
   U14924 : OAI22_X1 port map( A1 => n104_port, A2 => n11590, B1 => n232_port, 
                           B2 => n11573, ZN => n7751);
   U14925 : AOI21_X1 port map( B1 => n7766, B2 => n7767, A => n11069, ZN => 
                           n7765);
   U14926 : AOI221_X1 port map( B1 => n11015, B2 => n10337, C1 => n10998, C2 =>
                           n9889, A => n7769, ZN => n7766);
   U14927 : AOI221_X1 port map( B1 => n11051, B2 => n10338, C1 => n11033, C2 =>
                           n9890, A => n7768, ZN => n7767);
   U14928 : OAI22_X1 port map( A1 => n103_port, A2 => n11590, B1 => n231_port, 
                           B2 => n11573, ZN => n7769);
   U14929 : AOI21_X1 port map( B1 => n7784, B2 => n7785, A => n11069, ZN => 
                           n7783);
   U14930 : AOI221_X1 port map( B1 => n11016, B2 => n10339, C1 => n10999, C2 =>
                           n9891, A => n7787, ZN => n7784);
   U14931 : AOI221_X1 port map( B1 => n11051, B2 => n10340, C1 => n11033, C2 =>
                           n9892, A => n7786, ZN => n7785);
   U14932 : OAI22_X1 port map( A1 => n102_port, A2 => n11590, B1 => n230_port, 
                           B2 => n11573, ZN => n7787);
   U14933 : AOI21_X1 port map( B1 => n7802, B2 => n7803, A => n11069, ZN => 
                           n7801);
   U14934 : AOI221_X1 port map( B1 => n11016, B2 => n10341, C1 => n10999, C2 =>
                           n9893, A => n7805, ZN => n7802);
   U14935 : AOI221_X1 port map( B1 => n11051, B2 => n10342, C1 => n11033, C2 =>
                           n9894, A => n7804, ZN => n7803);
   U14936 : OAI22_X1 port map( A1 => n101_port, A2 => n11590, B1 => n229_port, 
                           B2 => n11573, ZN => n7805);
   U14937 : AOI21_X1 port map( B1 => n7820, B2 => n7821, A => n11068, ZN => 
                           n7819);
   U14938 : AOI221_X1 port map( B1 => n11016, B2 => n10343, C1 => n10999, C2 =>
                           n9895, A => n7823, ZN => n7820);
   U14939 : AOI221_X1 port map( B1 => n11051, B2 => n10344, C1 => n11033, C2 =>
                           n9896, A => n7822, ZN => n7821);
   U14940 : OAI22_X1 port map( A1 => n100_port, A2 => n11589, B1 => n228_port, 
                           B2 => n11572, ZN => n7823);
   U14941 : AOI21_X1 port map( B1 => n7838, B2 => n7839, A => n11068, ZN => 
                           n7837);
   U14942 : AOI221_X1 port map( B1 => n11016, B2 => n10345, C1 => n10999, C2 =>
                           n9897, A => n7841, ZN => n7838);
   U14943 : AOI221_X1 port map( B1 => n11051, B2 => n10346, C1 => n11033, C2 =>
                           n9898, A => n7840, ZN => n7839);
   U14944 : OAI22_X1 port map( A1 => n99_port, A2 => n11589, B1 => n227_port, 
                           B2 => n11572, ZN => n7841);
   U14945 : AOI21_X1 port map( B1 => n7856, B2 => n7857, A => n11068, ZN => 
                           n7855);
   U14946 : AOI221_X1 port map( B1 => n11016, B2 => n10347, C1 => n10999, C2 =>
                           n9899, A => n7859, ZN => n7856);
   U14947 : AOI221_X1 port map( B1 => n11051, B2 => n10348, C1 => n11034, C2 =>
                           n9900, A => n7858, ZN => n7857);
   U14948 : OAI22_X1 port map( A1 => n98_port, A2 => n11589, B1 => n226_port, 
                           B2 => n11572, ZN => n7859);
   U14949 : AOI21_X1 port map( B1 => n7874, B2 => n7875, A => n11068, ZN => 
                           n7873);
   U14950 : AOI221_X1 port map( B1 => n11016, B2 => n10349, C1 => n10999, C2 =>
                           n9901, A => n7877, ZN => n7874);
   U14951 : AOI221_X1 port map( B1 => n11052, B2 => n10350, C1 => n11034, C2 =>
                           n9902, A => n7876, ZN => n7875);
   U14952 : OAI22_X1 port map( A1 => n97_port, A2 => n11589, B1 => n225_port, 
                           B2 => n11572, ZN => n7877);
   U14953 : AOI21_X1 port map( B1 => n7892, B2 => n7893, A => n11068, ZN => 
                           n7891);
   U14954 : AOI221_X1 port map( B1 => n11016, B2 => n10351, C1 => n10999, C2 =>
                           n9903, A => n7895, ZN => n7892);
   U14955 : AOI221_X1 port map( B1 => n11052, B2 => n10352, C1 => n11034, C2 =>
                           n9904, A => n7894, ZN => n7893);
   U14956 : OAI22_X1 port map( A1 => n96_port, A2 => n11589, B1 => n224_port, 
                           B2 => n11572, ZN => n7895);
   U14957 : AOI21_X1 port map( B1 => n7910, B2 => n7911, A => n11068, ZN => 
                           n7909);
   U14958 : AOI221_X1 port map( B1 => n11017, B2 => n10353, C1 => n11000, C2 =>
                           n9905, A => n7913, ZN => n7910);
   U14959 : AOI221_X1 port map( B1 => n11052, B2 => n10354, C1 => n11034, C2 =>
                           n9906, A => n7912, ZN => n7911);
   U14960 : OAI22_X1 port map( A1 => n95_port, A2 => n11589, B1 => n223_port, 
                           B2 => n11572, ZN => n7913);
   U14961 : AOI21_X1 port map( B1 => n7928, B2 => n7929, A => n11068, ZN => 
                           n7927);
   U14962 : AOI221_X1 port map( B1 => n11017, B2 => n10355, C1 => n11000, C2 =>
                           n9907, A => n7931, ZN => n7928);
   U14963 : AOI221_X1 port map( B1 => n11052, B2 => n10356, C1 => n11034, C2 =>
                           n9908, A => n7930, ZN => n7929);
   U14964 : OAI22_X1 port map( A1 => n94_port, A2 => n11588, B1 => n222_port, 
                           B2 => n11571, ZN => n7931);
   U14965 : AOI21_X1 port map( B1 => n7946, B2 => n7947, A => n11068, ZN => 
                           n7945);
   U14966 : AOI221_X1 port map( B1 => n11017, B2 => n10357, C1 => n11000, C2 =>
                           n9909, A => n7949, ZN => n7946);
   U14967 : AOI221_X1 port map( B1 => n11052, B2 => n10358, C1 => n11034, C2 =>
                           n9910, A => n7948, ZN => n7947);
   U14968 : OAI22_X1 port map( A1 => n93_port, A2 => n11588, B1 => n221_port, 
                           B2 => n11571, ZN => n7949);
   U14969 : AOI21_X1 port map( B1 => n7964, B2 => n7965, A => n11068, ZN => 
                           n7963);
   U14970 : AOI221_X1 port map( B1 => n11017, B2 => n10359, C1 => n11000, C2 =>
                           n9911, A => n7967, ZN => n7964);
   U14971 : AOI221_X1 port map( B1 => n11053, B2 => n10360, C1 => n11035, C2 =>
                           n9912, A => n7966, ZN => n7965);
   U14972 : OAI22_X1 port map( A1 => n92_port, A2 => n11588, B1 => n220_port, 
                           B2 => n11571, ZN => n7967);
   U14973 : AOI21_X1 port map( B1 => n7982, B2 => n7983, A => n11068, ZN => 
                           n7981);
   U14974 : AOI221_X1 port map( B1 => n11017, B2 => n10361, C1 => n11000, C2 =>
                           n9913, A => n7985, ZN => n7982);
   U14975 : AOI221_X1 port map( B1 => n11053, B2 => n10362, C1 => n11035, C2 =>
                           n9914, A => n7984, ZN => n7983);
   U14976 : OAI22_X1 port map( A1 => n91_port, A2 => n11588, B1 => n219_port, 
                           B2 => n11571, ZN => n7985);
   U14977 : AOI21_X1 port map( B1 => n8000, B2 => n8001, A => n11068, ZN => 
                           n7999);
   U14978 : AOI221_X1 port map( B1 => n11017, B2 => n10363, C1 => n11000, C2 =>
                           n9915, A => n8003, ZN => n8000);
   U14979 : AOI221_X1 port map( B1 => n11053, B2 => n10364, C1 => n11035, C2 =>
                           n9916, A => n8002, ZN => n8001);
   U14980 : OAI22_X1 port map( A1 => n90_port, A2 => n11588, B1 => n218_port, 
                           B2 => n11571, ZN => n8003);
   U14981 : AOI21_X1 port map( B1 => n8018, B2 => n8019, A => n11068, ZN => 
                           n8017);
   U14982 : AOI221_X1 port map( B1 => n11018, B2 => n10365, C1 => n11001, C2 =>
                           n9917, A => n8021, ZN => n8018);
   U14983 : AOI221_X1 port map( B1 => n11053, B2 => n10366, C1 => n11035, C2 =>
                           n9918, A => n8020, ZN => n8019);
   U14984 : OAI22_X1 port map( A1 => n89_port, A2 => n11588, B1 => n217_port, 
                           B2 => n11571, ZN => n8021);
   U14985 : AOI21_X1 port map( B1 => n8036, B2 => n8037, A => n11067, ZN => 
                           n8035);
   U14986 : AOI221_X1 port map( B1 => n11018, B2 => n10367, C1 => n11001, C2 =>
                           n9919, A => n8039, ZN => n8036);
   U14987 : AOI221_X1 port map( B1 => n11053, B2 => n10368, C1 => n11035, C2 =>
                           n9920, A => n8038, ZN => n8037);
   U14988 : OAI22_X1 port map( A1 => n88_port, A2 => n11587, B1 => n216_port, 
                           B2 => n11570, ZN => n8039);
   U14989 : AOI21_X1 port map( B1 => n8054, B2 => n8055, A => n11067, ZN => 
                           n8053);
   U14990 : AOI221_X1 port map( B1 => n11018, B2 => n10369, C1 => n11001, C2 =>
                           n9921, A => n8057, ZN => n8054);
   U14991 : AOI221_X1 port map( B1 => n11053, B2 => n10370, C1 => n11035, C2 =>
                           n9922, A => n8056, ZN => n8055);
   U14992 : OAI22_X1 port map( A1 => n87_port, A2 => n11587, B1 => n215_port, 
                           B2 => n11570, ZN => n8057);
   U14993 : AOI21_X1 port map( B1 => n8072, B2 => n8073, A => n11067, ZN => 
                           n8071);
   U14994 : AOI221_X1 port map( B1 => n11018, B2 => n10371, C1 => n11001, C2 =>
                           n9923, A => n8075, ZN => n8072);
   U14995 : AOI221_X1 port map( B1 => n11054, B2 => n10372, C1 => n11036, C2 =>
                           n9924, A => n8074, ZN => n8073);
   U14996 : OAI22_X1 port map( A1 => n86_port, A2 => n11587, B1 => n214_port, 
                           B2 => n11570, ZN => n8075);
   U14997 : AOI21_X1 port map( B1 => n8090, B2 => n8091, A => n11067, ZN => 
                           n8089);
   U14998 : AOI221_X1 port map( B1 => n11018, B2 => n10373, C1 => n11001, C2 =>
                           n9925, A => n8093, ZN => n8090);
   U14999 : AOI221_X1 port map( B1 => n11054, B2 => n10374, C1 => n11036, C2 =>
                           n9926, A => n8092, ZN => n8091);
   U15000 : OAI22_X1 port map( A1 => n85_port, A2 => n11587, B1 => n213_port, 
                           B2 => n11570, ZN => n8093);
   U15001 : AOI21_X1 port map( B1 => n8108, B2 => n8109, A => n11067, ZN => 
                           n8107);
   U15002 : AOI221_X1 port map( B1 => n11018, B2 => n10375, C1 => n11001, C2 =>
                           n9927, A => n8111, ZN => n8108);
   U15003 : AOI221_X1 port map( B1 => n11054, B2 => n10376, C1 => n11036, C2 =>
                           n9928, A => n8110, ZN => n8109);
   U15004 : OAI22_X1 port map( A1 => n84_port, A2 => n11587, B1 => n212_port, 
                           B2 => n11570, ZN => n8111);
   U15005 : AOI21_X1 port map( B1 => n8126, B2 => n8127, A => n11067, ZN => 
                           n8125);
   U15006 : AOI221_X1 port map( B1 => n11019, B2 => n10377, C1 => n11002, C2 =>
                           n9929, A => n8129, ZN => n8126);
   U15007 : AOI221_X1 port map( B1 => n11054, B2 => n10378, C1 => n11036, C2 =>
                           n9930, A => n8128, ZN => n8127);
   U15008 : OAI22_X1 port map( A1 => n83_port, A2 => n11587, B1 => n211_port, 
                           B2 => n11570, ZN => n8129);
   U15009 : AOI21_X1 port map( B1 => n8144, B2 => n8145, A => n11067, ZN => 
                           n8143);
   U15010 : AOI221_X1 port map( B1 => n11019, B2 => n10379, C1 => n11002, C2 =>
                           n9931, A => n8147, ZN => n8144);
   U15011 : AOI221_X1 port map( B1 => n11054, B2 => n10380, C1 => n11036, C2 =>
                           n9932, A => n8146, ZN => n8145);
   U15012 : OAI22_X1 port map( A1 => n82_port, A2 => n11586, B1 => n210_port, 
                           B2 => n11569, ZN => n8147);
   U15013 : AOI21_X1 port map( B1 => n8162, B2 => n8163, A => n11067, ZN => 
                           n8161);
   U15014 : AOI221_X1 port map( B1 => n11019, B2 => n10381, C1 => n11002, C2 =>
                           n9933, A => n8165, ZN => n8162);
   U15015 : AOI221_X1 port map( B1 => n11054, B2 => n10382, C1 => n11036, C2 =>
                           n9934, A => n8164, ZN => n8163);
   U15016 : OAI22_X1 port map( A1 => n81_port, A2 => n11586, B1 => n209_port, 
                           B2 => n11569, ZN => n8165);
   U15017 : AOI21_X1 port map( B1 => n8180, B2 => n8181, A => n11067, ZN => 
                           n8179);
   U15018 : AOI221_X1 port map( B1 => n11019, B2 => n10383, C1 => n11002, C2 =>
                           n9935, A => n8183, ZN => n8180);
   U15019 : AOI221_X1 port map( B1 => n11055, B2 => n10384, C1 => n11037, C2 =>
                           n9936, A => n8182, ZN => n8181);
   U15020 : OAI22_X1 port map( A1 => n80_port, A2 => n11586, B1 => n208_port, 
                           B2 => n11569, ZN => n8183);
   U15021 : AOI21_X1 port map( B1 => n8198, B2 => n8199, A => n11067, ZN => 
                           n8197);
   U15022 : AOI221_X1 port map( B1 => n11019, B2 => n10385, C1 => n11002, C2 =>
                           n9937, A => n8201, ZN => n8198);
   U15023 : AOI221_X1 port map( B1 => n11055, B2 => n10386, C1 => n11037, C2 =>
                           n9938, A => n8200, ZN => n8199);
   U15024 : OAI22_X1 port map( A1 => n79_port, A2 => n11586, B1 => n207_port, 
                           B2 => n11569, ZN => n8201);
   U15025 : AOI21_X1 port map( B1 => n8216, B2 => n8217, A => n11067, ZN => 
                           n8215);
   U15026 : AOI221_X1 port map( B1 => n11019, B2 => n10387, C1 => n11002, C2 =>
                           n9939, A => n8219, ZN => n8216);
   U15027 : AOI221_X1 port map( B1 => n11055, B2 => n10388, C1 => n11037, C2 =>
                           n9940, A => n8218, ZN => n8217);
   U15028 : OAI22_X1 port map( A1 => n78_port, A2 => n11586, B1 => n206_port, 
                           B2 => n11569, ZN => n8219);
   U15029 : AOI21_X1 port map( B1 => n8234, B2 => n8235, A => n11067, ZN => 
                           n8233);
   U15030 : AOI221_X1 port map( B1 => n11019, B2 => n10389, C1 => n11002, C2 =>
                           n9941, A => n8237, ZN => n8234);
   U15031 : AOI221_X1 port map( B1 => n11055, B2 => n10390, C1 => n11037, C2 =>
                           n9942, A => n8236, ZN => n8235);
   U15032 : OAI22_X1 port map( A1 => n77_port, A2 => n11586, B1 => n205_port, 
                           B2 => n11569, ZN => n8237);
   U15033 : AOI21_X1 port map( B1 => n8252, B2 => n8253, A => n11066, ZN => 
                           n8251);
   U15034 : AOI221_X1 port map( B1 => n11020, B2 => n10391, C1 => n11003, C2 =>
                           n9943, A => n8255, ZN => n8252);
   U15035 : AOI221_X1 port map( B1 => n11055, B2 => n10392, C1 => n11037, C2 =>
                           n9944, A => n8254, ZN => n8253);
   U15036 : OAI22_X1 port map( A1 => n76_port, A2 => n11585, B1 => n204_port, 
                           B2 => n11568, ZN => n8255);
   U15037 : AOI21_X1 port map( B1 => n8270, B2 => n8271, A => n11066, ZN => 
                           n8269);
   U15038 : AOI221_X1 port map( B1 => n11020, B2 => n10393, C1 => n11003, C2 =>
                           n9945, A => n8273, ZN => n8270);
   U15039 : AOI221_X1 port map( B1 => n11055, B2 => n10394, C1 => n11037, C2 =>
                           n9946, A => n8272, ZN => n8271);
   U15040 : OAI22_X1 port map( A1 => n75_port, A2 => n11585, B1 => n203_port, 
                           B2 => n11568, ZN => n8273);
   U15041 : AOI21_X1 port map( B1 => n8288, B2 => n8289, A => n11066, ZN => 
                           n8287);
   U15042 : AOI221_X1 port map( B1 => n11020, B2 => n10395, C1 => n11003, C2 =>
                           n9947, A => n8291, ZN => n8288);
   U15043 : AOI221_X1 port map( B1 => n11056, B2 => n10396, C1 => n11038, C2 =>
                           n9948, A => n8290, ZN => n8289);
   U15044 : OAI22_X1 port map( A1 => n74_port, A2 => n11585, B1 => n202_port, 
                           B2 => n11568, ZN => n8291);
   U15045 : AOI21_X1 port map( B1 => n8306, B2 => n8307, A => n11066, ZN => 
                           n8305);
   U15046 : AOI221_X1 port map( B1 => n11020, B2 => n10397, C1 => n11003, C2 =>
                           n9949, A => n8309, ZN => n8306);
   U15047 : AOI221_X1 port map( B1 => n11056, B2 => n10398, C1 => n11038, C2 =>
                           n9950, A => n8308, ZN => n8307);
   U15048 : OAI22_X1 port map( A1 => n73_port, A2 => n11585, B1 => n201_port, 
                           B2 => n11568, ZN => n8309);
   U15049 : AOI21_X1 port map( B1 => n8324, B2 => n8325, A => n11066, ZN => 
                           n8323);
   U15050 : AOI221_X1 port map( B1 => n11020, B2 => n10399, C1 => n11003, C2 =>
                           n9951, A => n8327, ZN => n8324);
   U15051 : AOI221_X1 port map( B1 => n11056, B2 => n10400, C1 => n11038, C2 =>
                           n9952, A => n8326, ZN => n8325);
   U15052 : OAI22_X1 port map( A1 => n72_port, A2 => n11585, B1 => n200_port, 
                           B2 => n11568, ZN => n8327);
   U15053 : AOI21_X1 port map( B1 => n8342, B2 => n8343, A => n11066, ZN => 
                           n8341);
   U15054 : AOI221_X1 port map( B1 => n11020, B2 => n10401, C1 => n11003, C2 =>
                           n9953, A => n8345, ZN => n8342);
   U15055 : AOI221_X1 port map( B1 => n11056, B2 => n10402, C1 => n11038, C2 =>
                           n9954, A => n8344, ZN => n8343);
   U15056 : OAI22_X1 port map( A1 => n71_port, A2 => n11585, B1 => n199_port, 
                           B2 => n11568, ZN => n8345);
   U15057 : AOI21_X1 port map( B1 => n8360, B2 => n8361, A => n11066, ZN => 
                           n8359);
   U15058 : AOI221_X1 port map( B1 => n11021, B2 => n10403, C1 => n11004, C2 =>
                           n9955, A => n8363, ZN => n8360);
   U15059 : AOI221_X1 port map( B1 => n11056, B2 => n10404, C1 => n11038, C2 =>
                           n9956, A => n8362, ZN => n8361);
   U15060 : OAI22_X1 port map( A1 => n70_port, A2 => n11584, B1 => n198_port, 
                           B2 => n11567, ZN => n8363);
   U15061 : AOI21_X1 port map( B1 => n8378, B2 => n8379, A => n11066, ZN => 
                           n8377);
   U15062 : AOI221_X1 port map( B1 => n11021, B2 => n10405, C1 => n11004, C2 =>
                           n9957, A => n8381, ZN => n8378);
   U15063 : AOI221_X1 port map( B1 => n11056, B2 => n10406, C1 => n11038, C2 =>
                           n9958, A => n8380, ZN => n8379);
   U15064 : OAI22_X1 port map( A1 => n69_port, A2 => n11584, B1 => n197_port, 
                           B2 => n11567, ZN => n8381);
   U15065 : AOI21_X1 port map( B1 => n8396, B2 => n8397, A => n11066, ZN => 
                           n8395);
   U15066 : AOI221_X1 port map( B1 => n11021, B2 => n10407, C1 => n11004, C2 =>
                           n9959, A => n8399, ZN => n8396);
   U15067 : AOI221_X1 port map( B1 => n11057, B2 => n10408, C1 => n11039, C2 =>
                           n9960, A => n8398, ZN => n8397);
   U15068 : OAI22_X1 port map( A1 => n68_port, A2 => n11584, B1 => n196_port, 
                           B2 => n11567, ZN => n8399);
   U15069 : AOI21_X1 port map( B1 => n8414, B2 => n8415, A => n11066, ZN => 
                           n8413);
   U15070 : AOI221_X1 port map( B1 => n11021, B2 => n10409, C1 => n11004, C2 =>
                           n9961, A => n8417, ZN => n8414);
   U15071 : AOI221_X1 port map( B1 => n11057, B2 => n10410, C1 => n11039, C2 =>
                           n9962, A => n8416, ZN => n8415);
   U15072 : OAI22_X1 port map( A1 => n67_port, A2 => n11584, B1 => n195_port, 
                           B2 => n11567, ZN => n8417);
   U15073 : AOI21_X1 port map( B1 => n8432, B2 => n8433, A => n11066, ZN => 
                           n8431);
   U15074 : AOI221_X1 port map( B1 => n11021, B2 => n10411, C1 => n11004, C2 =>
                           n9963, A => n8435, ZN => n8432);
   U15075 : AOI221_X1 port map( B1 => n11057, B2 => n10412, C1 => n11039, C2 =>
                           n9964, A => n8434, ZN => n8433);
   U15076 : OAI22_X1 port map( A1 => n66_port, A2 => n11584, B1 => n194_port, 
                           B2 => n11567, ZN => n8435);
   U15077 : AOI21_X1 port map( B1 => n8450, B2 => n8451, A => n11066, ZN => 
                           n8449);
   U15078 : AOI221_X1 port map( B1 => n11021, B2 => n10413, C1 => n11004, C2 =>
                           n9965, A => n8453, ZN => n8450);
   U15079 : AOI221_X1 port map( B1 => n11057, B2 => n10414, C1 => n11039, C2 =>
                           n9966, A => n8452, ZN => n8451);
   U15080 : OAI22_X1 port map( A1 => n65_port, A2 => n11584, B1 => n193_port, 
                           B2 => n11567, ZN => n8453);
   U15081 : AOI21_X1 port map( B1 => n8474, B2 => n8475, A => n10846, ZN => 
                           n8473);
   U15082 : AOI221_X1 port map( B1 => n10792, B2 => n10287, C1 => n10775, C2 =>
                           n9839, A => n8482, ZN => n8474);
   U15083 : AOI221_X1 port map( B1 => n10827, B2 => n10288, C1 => n10804, C2 =>
                           n9840, A => n8479, ZN => n8475);
   U15084 : OAI22_X1 port map( A1 => n128_port, A2 => n11662, B1 => n256_port, 
                           B2 => n11645, ZN => n8482);
   U15085 : AOI21_X1 port map( B1 => n8514, B2 => n8515, A => n10846, ZN => 
                           n8513);
   U15086 : AOI221_X1 port map( B1 => n10787, B2 => n10289, C1 => n10770, C2 =>
                           n9841, A => n8517, ZN => n8514);
   U15087 : AOI221_X1 port map( B1 => n10822, B2 => n10290, C1 => n10804, C2 =>
                           n9842, A => n8516, ZN => n8515);
   U15088 : OAI22_X1 port map( A1 => n127_port, A2 => n11662, B1 => n255_port, 
                           B2 => n11645, ZN => n8517);
   U15089 : AOI21_X1 port map( B1 => n8532, B2 => n8533, A => n10846, ZN => 
                           n8531);
   U15090 : AOI221_X1 port map( B1 => n10787, B2 => n10291, C1 => n10770, C2 =>
                           n9843, A => n8535, ZN => n8532);
   U15091 : AOI221_X1 port map( B1 => n10822, B2 => n10292, C1 => n10804, C2 =>
                           n9844, A => n8534, ZN => n8533);
   U15092 : OAI22_X1 port map( A1 => n126_port, A2 => n11662, B1 => n254_port, 
                           B2 => n11645, ZN => n8535);
   U15093 : AOI21_X1 port map( B1 => n8550, B2 => n8551, A => n10846, ZN => 
                           n8549);
   U15094 : AOI221_X1 port map( B1 => n10787, B2 => n10293, C1 => n10770, C2 =>
                           n9845, A => n8553, ZN => n8550);
   U15095 : AOI221_X1 port map( B1 => n10822, B2 => n10294, C1 => n10804, C2 =>
                           n9846, A => n8552, ZN => n8551);
   U15096 : OAI22_X1 port map( A1 => n125_port, A2 => n11662, B1 => n253_port, 
                           B2 => n11645, ZN => n8553);
   U15097 : AOI21_X1 port map( B1 => n8568, B2 => n8569, A => n10845, ZN => 
                           n8567);
   U15098 : AOI221_X1 port map( B1 => n10787, B2 => n10295, C1 => n10770, C2 =>
                           n9847, A => n8571, ZN => n8568);
   U15099 : AOI221_X1 port map( B1 => n10822, B2 => n10296, C1 => n10804, C2 =>
                           n9848, A => n8570, ZN => n8569);
   U15100 : OAI22_X1 port map( A1 => n124_port, A2 => n11661, B1 => n252_port, 
                           B2 => n11644, ZN => n8571);
   U15101 : AOI21_X1 port map( B1 => n8586, B2 => n8587, A => n10845, ZN => 
                           n8585);
   U15102 : AOI221_X1 port map( B1 => n10787, B2 => n10297, C1 => n10770, C2 =>
                           n9849, A => n8589, ZN => n8586);
   U15103 : AOI221_X1 port map( B1 => n10822, B2 => n10298, C1 => n10804, C2 =>
                           n9850, A => n8588, ZN => n8587);
   U15104 : OAI22_X1 port map( A1 => n123_port, A2 => n11661, B1 => n251_port, 
                           B2 => n11644, ZN => n8589);
   U15105 : AOI21_X1 port map( B1 => n8604, B2 => n8605, A => n10845, ZN => 
                           n8603);
   U15106 : AOI221_X1 port map( B1 => n10787, B2 => n10299, C1 => n10770, C2 =>
                           n9851, A => n8607, ZN => n8604);
   U15107 : AOI221_X1 port map( B1 => n10822, B2 => n10300, C1 => n10805, C2 =>
                           n9852, A => n8606, ZN => n8605);
   U15108 : OAI22_X1 port map( A1 => n122_port, A2 => n11661, B1 => n250_port, 
                           B2 => n11644, ZN => n8607);
   U15109 : AOI21_X1 port map( B1 => n8622, B2 => n8623, A => n10845, ZN => 
                           n8621);
   U15110 : AOI221_X1 port map( B1 => n10788, B2 => n10301, C1 => n10771, C2 =>
                           n9853, A => n8625, ZN => n8622);
   U15111 : AOI221_X1 port map( B1 => n10823, B2 => n10302, C1 => n10805, C2 =>
                           n9854, A => n8624, ZN => n8623);
   U15112 : OAI22_X1 port map( A1 => n121_port, A2 => n11661, B1 => n249_port, 
                           B2 => n11644, ZN => n8625);
   U15113 : AOI21_X1 port map( B1 => n8640, B2 => n8641, A => n10845, ZN => 
                           n8639);
   U15114 : AOI221_X1 port map( B1 => n10788, B2 => n10303, C1 => n10771, C2 =>
                           n9855, A => n8643, ZN => n8640);
   U15115 : AOI221_X1 port map( B1 => n10823, B2 => n10304, C1 => n10805, C2 =>
                           n9856, A => n8642, ZN => n8641);
   U15116 : OAI22_X1 port map( A1 => n120_port, A2 => n11661, B1 => n248_port, 
                           B2 => n11644, ZN => n8643);
   U15117 : AOI21_X1 port map( B1 => n8658, B2 => n8659, A => n10845, ZN => 
                           n8657);
   U15118 : AOI221_X1 port map( B1 => n10788, B2 => n10305, C1 => n10771, C2 =>
                           n9857, A => n8661, ZN => n8658);
   U15119 : AOI221_X1 port map( B1 => n10823, B2 => n10306, C1 => n10805, C2 =>
                           n9858, A => n8660, ZN => n8659);
   U15120 : OAI22_X1 port map( A1 => n119_port, A2 => n11661, B1 => n247_port, 
                           B2 => n11644, ZN => n8661);
   U15121 : AOI21_X1 port map( B1 => n8676, B2 => n8677, A => n10845, ZN => 
                           n8675);
   U15122 : AOI221_X1 port map( B1 => n10788, B2 => n10307, C1 => n10771, C2 =>
                           n9859, A => n8679, ZN => n8676);
   U15123 : AOI221_X1 port map( B1 => n10823, B2 => n10308, C1 => n10805, C2 =>
                           n9860, A => n8678, ZN => n8677);
   U15124 : OAI22_X1 port map( A1 => n118_port, A2 => n11660, B1 => n246_port, 
                           B2 => n11643, ZN => n8679);
   U15125 : AOI21_X1 port map( B1 => n8694, B2 => n8695, A => n10845, ZN => 
                           n8693);
   U15126 : AOI221_X1 port map( B1 => n10788, B2 => n10309, C1 => n10771, C2 =>
                           n9861, A => n8697, ZN => n8694);
   U15127 : AOI221_X1 port map( B1 => n10823, B2 => n10310, C1 => n10805, C2 =>
                           n9862, A => n8696, ZN => n8695);
   U15128 : OAI22_X1 port map( A1 => n117_port, A2 => n11660, B1 => n245_port, 
                           B2 => n11643, ZN => n8697);
   U15129 : AOI21_X1 port map( B1 => n8712, B2 => n8713, A => n10845, ZN => 
                           n8711);
   U15130 : AOI221_X1 port map( B1 => n10788, B2 => n10311, C1 => n10771, C2 =>
                           n9863, A => n8715, ZN => n8712);
   U15131 : AOI221_X1 port map( B1 => n10823, B2 => n10312, C1 => n10806, C2 =>
                           n9864, A => n8714, ZN => n8713);
   U15132 : OAI22_X1 port map( A1 => n116_port, A2 => n11660, B1 => n244_port, 
                           B2 => n11643, ZN => n8715);
   U15133 : AOI21_X1 port map( B1 => n8730, B2 => n8731, A => n10845, ZN => 
                           n8729);
   U15134 : AOI221_X1 port map( B1 => n10789, B2 => n10313, C1 => n10772, C2 =>
                           n9865, A => n8733, ZN => n8730);
   U15135 : AOI221_X1 port map( B1 => n10824, B2 => n10314, C1 => n10806, C2 =>
                           n9866, A => n8732, ZN => n8731);
   U15136 : OAI22_X1 port map( A1 => n115_port, A2 => n11660, B1 => n243_port, 
                           B2 => n11643, ZN => n8733);
   U15137 : AOI21_X1 port map( B1 => n8748, B2 => n8749, A => n10845, ZN => 
                           n8747);
   U15138 : AOI221_X1 port map( B1 => n10789, B2 => n10315, C1 => n10772, C2 =>
                           n9867, A => n8751, ZN => n8748);
   U15139 : AOI221_X1 port map( B1 => n10824, B2 => n10316, C1 => n10806, C2 =>
                           n9868, A => n8750, ZN => n8749);
   U15140 : OAI22_X1 port map( A1 => n114_port, A2 => n11660, B1 => n242_port, 
                           B2 => n11643, ZN => n8751);
   U15141 : AOI21_X1 port map( B1 => n8766, B2 => n8767, A => n10845, ZN => 
                           n8765);
   U15142 : AOI221_X1 port map( B1 => n10789, B2 => n10317, C1 => n10772, C2 =>
                           n9869, A => n8769, ZN => n8766);
   U15143 : AOI221_X1 port map( B1 => n10824, B2 => n10318, C1 => n10806, C2 =>
                           n9870, A => n8768, ZN => n8767);
   U15144 : OAI22_X1 port map( A1 => n113_port, A2 => n11660, B1 => n241_port, 
                           B2 => n11643, ZN => n8769);
   U15145 : AOI21_X1 port map( B1 => n8784, B2 => n8785, A => n10844, ZN => 
                           n8783);
   U15146 : AOI221_X1 port map( B1 => n10789, B2 => n10319, C1 => n10772, C2 =>
                           n9871, A => n8787, ZN => n8784);
   U15147 : AOI221_X1 port map( B1 => n10824, B2 => n10320, C1 => n10806, C2 =>
                           n9872, A => n8786, ZN => n8785);
   U15148 : OAI22_X1 port map( A1 => n112_port, A2 => n11659, B1 => n240_port, 
                           B2 => n11642, ZN => n8787);
   U15149 : AOI21_X1 port map( B1 => n8802, B2 => n8803, A => n10844, ZN => 
                           n8801);
   U15150 : AOI221_X1 port map( B1 => n10789, B2 => n10321, C1 => n10772, C2 =>
                           n9873, A => n8805, ZN => n8802);
   U15151 : AOI221_X1 port map( B1 => n10824, B2 => n10322, C1 => n10806, C2 =>
                           n9874, A => n8804, ZN => n8803);
   U15152 : OAI22_X1 port map( A1 => n111_port, A2 => n11659, B1 => n239_port, 
                           B2 => n11642, ZN => n8805);
   U15153 : AOI21_X1 port map( B1 => n8820, B2 => n8821, A => n10844, ZN => 
                           n8819);
   U15154 : AOI221_X1 port map( B1 => n10789, B2 => n10323, C1 => n10772, C2 =>
                           n9875, A => n8823, ZN => n8820);
   U15155 : AOI221_X1 port map( B1 => n10824, B2 => n10324, C1 => n10807, C2 =>
                           n9876, A => n8822, ZN => n8821);
   U15156 : OAI22_X1 port map( A1 => n110_port, A2 => n11659, B1 => n238_port, 
                           B2 => n11642, ZN => n8823);
   U15157 : AOI21_X1 port map( B1 => n8838, B2 => n8839, A => n10844, ZN => 
                           n8837);
   U15158 : AOI221_X1 port map( B1 => n10789, B2 => n10325, C1 => n10772, C2 =>
                           n9877, A => n8841, ZN => n8838);
   U15159 : AOI221_X1 port map( B1 => n10825, B2 => n10326, C1 => n10807, C2 =>
                           n9878, A => n8840, ZN => n8839);
   U15160 : OAI22_X1 port map( A1 => n109_port, A2 => n11659, B1 => n237_port, 
                           B2 => n11642, ZN => n8841);
   U15161 : AOI21_X1 port map( B1 => n8856, B2 => n8857, A => n10844, ZN => 
                           n8855);
   U15162 : AOI221_X1 port map( B1 => n10790, B2 => n10327, C1 => n10773, C2 =>
                           n9879, A => n8859, ZN => n8856);
   U15163 : AOI221_X1 port map( B1 => n10825, B2 => n10328, C1 => n10807, C2 =>
                           n9880, A => n8858, ZN => n8857);
   U15164 : OAI22_X1 port map( A1 => n108_port, A2 => n11659, B1 => n236_port, 
                           B2 => n11642, ZN => n8859);
   U15165 : AOI21_X1 port map( B1 => n8874, B2 => n8875, A => n10844, ZN => 
                           n8873);
   U15166 : AOI221_X1 port map( B1 => n10790, B2 => n10329, C1 => n10773, C2 =>
                           n9881, A => n8877, ZN => n8874);
   U15167 : AOI221_X1 port map( B1 => n10825, B2 => n10330, C1 => n10807, C2 =>
                           n9882, A => n8876, ZN => n8875);
   U15168 : OAI22_X1 port map( A1 => n107_port, A2 => n11659, B1 => n235_port, 
                           B2 => n11642, ZN => n8877);
   U15169 : AOI21_X1 port map( B1 => n8892, B2 => n8893, A => n10844, ZN => 
                           n8891);
   U15170 : AOI221_X1 port map( B1 => n10790, B2 => n10331, C1 => n10773, C2 =>
                           n9883, A => n8895, ZN => n8892);
   U15171 : AOI221_X1 port map( B1 => n10825, B2 => n10332, C1 => n10807, C2 =>
                           n9884, A => n8894, ZN => n8893);
   U15172 : OAI22_X1 port map( A1 => n106_port, A2 => n11658, B1 => n234_port, 
                           B2 => n11641, ZN => n8895);
   U15173 : AOI21_X1 port map( B1 => n8910, B2 => n8911, A => n10844, ZN => 
                           n8909);
   U15174 : AOI221_X1 port map( B1 => n10790, B2 => n10333, C1 => n10773, C2 =>
                           n9885, A => n8913, ZN => n8910);
   U15175 : AOI221_X1 port map( B1 => n10825, B2 => n10334, C1 => n10807, C2 =>
                           n9886, A => n8912, ZN => n8911);
   U15176 : OAI22_X1 port map( A1 => n105_port, A2 => n11658, B1 => n233_port, 
                           B2 => n11641, ZN => n8913);
   U15177 : AOI21_X1 port map( B1 => n8928, B2 => n8929, A => n10844, ZN => 
                           n8927);
   U15178 : AOI221_X1 port map( B1 => n10790, B2 => n10335, C1 => n10773, C2 =>
                           n9887, A => n8931, ZN => n8928);
   U15179 : AOI221_X1 port map( B1 => n10825, B2 => n10336, C1 => n10808, C2 =>
                           n9888, A => n8930, ZN => n8929);
   U15180 : OAI22_X1 port map( A1 => n104_port, A2 => n11658, B1 => n232_port, 
                           B2 => n11641, ZN => n8931);
   U15181 : AOI21_X1 port map( B1 => n8946, B2 => n8947, A => n10844, ZN => 
                           n8945);
   U15182 : AOI221_X1 port map( B1 => n10790, B2 => n10337, C1 => n10773, C2 =>
                           n9889, A => n8949, ZN => n8946);
   U15183 : AOI221_X1 port map( B1 => n10826, B2 => n10338, C1 => n10808, C2 =>
                           n9890, A => n8948, ZN => n8947);
   U15184 : OAI22_X1 port map( A1 => n103_port, A2 => n11658, B1 => n231_port, 
                           B2 => n11641, ZN => n8949);
   U15185 : AOI21_X1 port map( B1 => n8964, B2 => n8965, A => n10844, ZN => 
                           n8963);
   U15186 : AOI221_X1 port map( B1 => n10791, B2 => n10339, C1 => n10774, C2 =>
                           n9891, A => n8967, ZN => n8964);
   U15187 : AOI221_X1 port map( B1 => n10826, B2 => n10340, C1 => n10808, C2 =>
                           n9892, A => n8966, ZN => n8965);
   U15188 : OAI22_X1 port map( A1 => n102_port, A2 => n11658, B1 => n230_port, 
                           B2 => n11641, ZN => n8967);
   U15189 : AOI21_X1 port map( B1 => n8982, B2 => n8983, A => n10844, ZN => 
                           n8981);
   U15190 : AOI221_X1 port map( B1 => n10791, B2 => n10341, C1 => n10774, C2 =>
                           n9893, A => n8985, ZN => n8982);
   U15191 : AOI221_X1 port map( B1 => n10826, B2 => n10342, C1 => n10808, C2 =>
                           n9894, A => n8984, ZN => n8983);
   U15192 : OAI22_X1 port map( A1 => n101_port, A2 => n11658, B1 => n229_port, 
                           B2 => n11641, ZN => n8985);
   U15193 : AOI21_X1 port map( B1 => n9000, B2 => n9001, A => n10843, ZN => 
                           n8999);
   U15194 : AOI221_X1 port map( B1 => n10791, B2 => n10343, C1 => n10774, C2 =>
                           n9895, A => n9003, ZN => n9000);
   U15195 : AOI221_X1 port map( B1 => n10826, B2 => n10344, C1 => n10808, C2 =>
                           n9896, A => n9002, ZN => n9001);
   U15196 : OAI22_X1 port map( A1 => n100_port, A2 => n11657, B1 => n228_port, 
                           B2 => n11640, ZN => n9003);
   U15197 : AOI21_X1 port map( B1 => n9018, B2 => n9019, A => n10843, ZN => 
                           n9017);
   U15198 : AOI221_X1 port map( B1 => n10791, B2 => n10345, C1 => n10774, C2 =>
                           n9897, A => n9021, ZN => n9018);
   U15199 : AOI221_X1 port map( B1 => n10826, B2 => n10346, C1 => n10808, C2 =>
                           n9898, A => n9020, ZN => n9019);
   U15200 : OAI22_X1 port map( A1 => n99_port, A2 => n11657, B1 => n227_port, 
                           B2 => n11640, ZN => n9021);
   U15201 : AOI21_X1 port map( B1 => n9036, B2 => n9037, A => n10843, ZN => 
                           n9035);
   U15202 : AOI221_X1 port map( B1 => n10791, B2 => n10347, C1 => n10774, C2 =>
                           n9899, A => n9039, ZN => n9036);
   U15203 : AOI221_X1 port map( B1 => n10826, B2 => n10348, C1 => n10809, C2 =>
                           n9900, A => n9038, ZN => n9037);
   U15204 : OAI22_X1 port map( A1 => n98_port, A2 => n11657, B1 => n226_port, 
                           B2 => n11640, ZN => n9039);
   U15205 : AOI21_X1 port map( B1 => n9054, B2 => n9055, A => n10843, ZN => 
                           n9053);
   U15206 : AOI221_X1 port map( B1 => n10791, B2 => n10349, C1 => n10774, C2 =>
                           n9901, A => n9057, ZN => n9054);
   U15207 : AOI221_X1 port map( B1 => n10827, B2 => n10350, C1 => n10809, C2 =>
                           n9902, A => n9056, ZN => n9055);
   U15208 : OAI22_X1 port map( A1 => n97_port, A2 => n11657, B1 => n225_port, 
                           B2 => n11640, ZN => n9057);
   U15209 : AOI21_X1 port map( B1 => n9072, B2 => n9073, A => n10843, ZN => 
                           n9071);
   U15210 : AOI221_X1 port map( B1 => n10791, B2 => n10351, C1 => n10774, C2 =>
                           n9903, A => n9075, ZN => n9072);
   U15211 : AOI221_X1 port map( B1 => n10827, B2 => n10352, C1 => n10809, C2 =>
                           n9904, A => n9074, ZN => n9073);
   U15212 : OAI22_X1 port map( A1 => n96_port, A2 => n11657, B1 => n224_port, 
                           B2 => n11640, ZN => n9075);
   U15213 : AOI21_X1 port map( B1 => n9090, B2 => n9091, A => n10843, ZN => 
                           n9089);
   U15214 : AOI221_X1 port map( B1 => n10792, B2 => n10353, C1 => n10775, C2 =>
                           n9905, A => n9093, ZN => n9090);
   U15215 : AOI221_X1 port map( B1 => n10827, B2 => n10354, C1 => n10809, C2 =>
                           n9906, A => n9092, ZN => n9091);
   U15216 : OAI22_X1 port map( A1 => n95_port, A2 => n11657, B1 => n223_port, 
                           B2 => n11640, ZN => n9093);
   U15217 : AOI21_X1 port map( B1 => n9108, B2 => n9109, A => n10843, ZN => 
                           n9107);
   U15218 : AOI221_X1 port map( B1 => n10792, B2 => n10355, C1 => n10775, C2 =>
                           n9907, A => n9111, ZN => n9108);
   U15219 : AOI221_X1 port map( B1 => n10827, B2 => n10356, C1 => n10809, C2 =>
                           n9908, A => n9110, ZN => n9109);
   U15220 : OAI22_X1 port map( A1 => n94_port, A2 => n11656, B1 => n222_port, 
                           B2 => n11639, ZN => n9111);
   U15221 : AOI21_X1 port map( B1 => n9126, B2 => n9127, A => n10843, ZN => 
                           n9125);
   U15222 : AOI221_X1 port map( B1 => n10792, B2 => n10357, C1 => n10775, C2 =>
                           n9909, A => n9129, ZN => n9126);
   U15223 : AOI221_X1 port map( B1 => n10827, B2 => n10358, C1 => n10809, C2 =>
                           n9910, A => n9128, ZN => n9127);
   U15224 : OAI22_X1 port map( A1 => n93_port, A2 => n11656, B1 => n221_port, 
                           B2 => n11639, ZN => n9129);
   U15225 : AOI21_X1 port map( B1 => n9144, B2 => n9145, A => n10843, ZN => 
                           n9143);
   U15226 : AOI221_X1 port map( B1 => n10792, B2 => n10359, C1 => n10775, C2 =>
                           n9911, A => n9147, ZN => n9144);
   U15227 : AOI221_X1 port map( B1 => n10828, B2 => n10360, C1 => n10810, C2 =>
                           n9912, A => n9146, ZN => n9145);
   U15228 : OAI22_X1 port map( A1 => n92_port, A2 => n11656, B1 => n220_port, 
                           B2 => n11639, ZN => n9147);
   U15229 : AOI21_X1 port map( B1 => n9162, B2 => n9163, A => n10843, ZN => 
                           n9161);
   U15230 : AOI221_X1 port map( B1 => n10792, B2 => n10361, C1 => n10775, C2 =>
                           n9913, A => n9165, ZN => n9162);
   U15231 : AOI221_X1 port map( B1 => n10828, B2 => n10362, C1 => n10810, C2 =>
                           n9914, A => n9164, ZN => n9163);
   U15232 : OAI22_X1 port map( A1 => n91_port, A2 => n11656, B1 => n219_port, 
                           B2 => n11639, ZN => n9165);
   U15233 : AOI21_X1 port map( B1 => n9180, B2 => n9181, A => n10843, ZN => 
                           n9179);
   U15234 : AOI221_X1 port map( B1 => n10792, B2 => n10363, C1 => n10775, C2 =>
                           n9915, A => n9183, ZN => n9180);
   U15235 : AOI221_X1 port map( B1 => n10828, B2 => n10364, C1 => n10810, C2 =>
                           n9916, A => n9182, ZN => n9181);
   U15236 : OAI22_X1 port map( A1 => n90_port, A2 => n11656, B1 => n218_port, 
                           B2 => n11639, ZN => n9183);
   U15237 : AOI21_X1 port map( B1 => n9198, B2 => n9199, A => n10843, ZN => 
                           n9197);
   U15238 : AOI221_X1 port map( B1 => n10793, B2 => n10365, C1 => n10776, C2 =>
                           n9917, A => n9201, ZN => n9198);
   U15239 : AOI221_X1 port map( B1 => n10828, B2 => n10366, C1 => n10810, C2 =>
                           n9918, A => n9200, ZN => n9199);
   U15240 : OAI22_X1 port map( A1 => n89_port, A2 => n11656, B1 => n217_port, 
                           B2 => n11639, ZN => n9201);
   U15241 : AOI21_X1 port map( B1 => n9216, B2 => n9217, A => n10842, ZN => 
                           n9215);
   U15242 : AOI221_X1 port map( B1 => n10793, B2 => n10367, C1 => n10776, C2 =>
                           n9919, A => n9219, ZN => n9216);
   U15243 : AOI221_X1 port map( B1 => n10828, B2 => n10368, C1 => n10810, C2 =>
                           n9920, A => n9218, ZN => n9217);
   U15244 : OAI22_X1 port map( A1 => n88_port, A2 => n11655, B1 => n216_port, 
                           B2 => n11638, ZN => n9219);
   U15245 : AOI21_X1 port map( B1 => n9234, B2 => n9235, A => n10842, ZN => 
                           n9233);
   U15246 : AOI221_X1 port map( B1 => n10793, B2 => n10369, C1 => n10776, C2 =>
                           n9921, A => n9237, ZN => n9234);
   U15247 : AOI221_X1 port map( B1 => n10828, B2 => n10370, C1 => n10810, C2 =>
                           n9922, A => n9236, ZN => n9235);
   U15248 : OAI22_X1 port map( A1 => n87_port, A2 => n11655, B1 => n215_port, 
                           B2 => n11638, ZN => n9237);
   U15249 : AOI21_X1 port map( B1 => n9252, B2 => n9253, A => n10842, ZN => 
                           n9251);
   U15250 : AOI221_X1 port map( B1 => n10793, B2 => n10371, C1 => n10776, C2 =>
                           n9923, A => n9255, ZN => n9252);
   U15251 : AOI221_X1 port map( B1 => n10829, B2 => n10372, C1 => n10811, C2 =>
                           n9924, A => n9254, ZN => n9253);
   U15252 : OAI22_X1 port map( A1 => n86_port, A2 => n11655, B1 => n214_port, 
                           B2 => n11638, ZN => n9255);
   U15253 : AOI21_X1 port map( B1 => n9270, B2 => n9271, A => n10842, ZN => 
                           n9269);
   U15254 : AOI221_X1 port map( B1 => n10793, B2 => n10373, C1 => n10776, C2 =>
                           n9925, A => n9273, ZN => n9270);
   U15255 : AOI221_X1 port map( B1 => n10829, B2 => n10374, C1 => n10811, C2 =>
                           n9926, A => n9272, ZN => n9271);
   U15256 : OAI22_X1 port map( A1 => n85_port, A2 => n11655, B1 => n213_port, 
                           B2 => n11638, ZN => n9273);
   U15257 : AOI21_X1 port map( B1 => n9288, B2 => n9289, A => n10842, ZN => 
                           n9287);
   U15258 : AOI221_X1 port map( B1 => n10793, B2 => n10375, C1 => n10776, C2 =>
                           n9927, A => n9291, ZN => n9288);
   U15259 : AOI221_X1 port map( B1 => n10829, B2 => n10376, C1 => n10811, C2 =>
                           n9928, A => n9290, ZN => n9289);
   U15260 : OAI22_X1 port map( A1 => n84_port, A2 => n11655, B1 => n212_port, 
                           B2 => n11638, ZN => n9291);
   U15261 : AOI21_X1 port map( B1 => n9306, B2 => n9307, A => n10842, ZN => 
                           n9305);
   U15262 : AOI221_X1 port map( B1 => n10794, B2 => n10377, C1 => n10777, C2 =>
                           n9929, A => n9309, ZN => n9306);
   U15263 : AOI221_X1 port map( B1 => n10829, B2 => n10378, C1 => n10811, C2 =>
                           n9930, A => n9308, ZN => n9307);
   U15264 : OAI22_X1 port map( A1 => n83_port, A2 => n11655, B1 => n211_port, 
                           B2 => n11638, ZN => n9309);
   U15265 : AOI21_X1 port map( B1 => n9324, B2 => n9325, A => n10842, ZN => 
                           n9323);
   U15266 : AOI221_X1 port map( B1 => n10794, B2 => n10379, C1 => n10777, C2 =>
                           n9931, A => n9327, ZN => n9324);
   U15267 : AOI221_X1 port map( B1 => n10829, B2 => n10380, C1 => n10811, C2 =>
                           n9932, A => n9326, ZN => n9325);
   U15268 : OAI22_X1 port map( A1 => n82_port, A2 => n11654, B1 => n210_port, 
                           B2 => n11637, ZN => n9327);
   U15269 : AOI21_X1 port map( B1 => n9342, B2 => n9343, A => n10842, ZN => 
                           n9341);
   U15270 : AOI221_X1 port map( B1 => n10794, B2 => n10381, C1 => n10777, C2 =>
                           n9933, A => n9345, ZN => n9342);
   U15271 : AOI221_X1 port map( B1 => n10829, B2 => n10382, C1 => n10811, C2 =>
                           n9934, A => n9344, ZN => n9343);
   U15272 : OAI22_X1 port map( A1 => n81_port, A2 => n11654, B1 => n209_port, 
                           B2 => n11637, ZN => n9345);
   U15273 : AOI21_X1 port map( B1 => n9360, B2 => n9361, A => n10842, ZN => 
                           n9359);
   U15274 : AOI221_X1 port map( B1 => n10794, B2 => n10383, C1 => n10777, C2 =>
                           n9935, A => n9363, ZN => n9360);
   U15275 : AOI221_X1 port map( B1 => n10830, B2 => n10384, C1 => n10812, C2 =>
                           n9936, A => n9362, ZN => n9361);
   U15276 : OAI22_X1 port map( A1 => n80_port, A2 => n11654, B1 => n208_port, 
                           B2 => n11637, ZN => n9363);
   U15277 : AOI21_X1 port map( B1 => n9378, B2 => n9379, A => n10842, ZN => 
                           n9377);
   U15278 : AOI221_X1 port map( B1 => n10794, B2 => n10385, C1 => n10777, C2 =>
                           n9937, A => n9381, ZN => n9378);
   U15279 : AOI221_X1 port map( B1 => n10830, B2 => n10386, C1 => n10812, C2 =>
                           n9938, A => n9380, ZN => n9379);
   U15280 : OAI22_X1 port map( A1 => n79_port, A2 => n11654, B1 => n207_port, 
                           B2 => n11637, ZN => n9381);
   U15281 : AOI21_X1 port map( B1 => n9396, B2 => n9397, A => n10842, ZN => 
                           n9395);
   U15282 : AOI221_X1 port map( B1 => n10794, B2 => n10387, C1 => n10777, C2 =>
                           n9939, A => n9399, ZN => n9396);
   U15283 : AOI221_X1 port map( B1 => n10830, B2 => n10388, C1 => n10812, C2 =>
                           n9940, A => n9398, ZN => n9397);
   U15284 : OAI22_X1 port map( A1 => n78_port, A2 => n11654, B1 => n206_port, 
                           B2 => n11637, ZN => n9399);
   U15285 : AOI21_X1 port map( B1 => n9414, B2 => n9415, A => n10842, ZN => 
                           n9413);
   U15286 : AOI221_X1 port map( B1 => n10794, B2 => n10389, C1 => n10777, C2 =>
                           n9941, A => n9417, ZN => n9414);
   U15287 : AOI221_X1 port map( B1 => n10830, B2 => n10390, C1 => n10812, C2 =>
                           n9942, A => n9416, ZN => n9415);
   U15288 : OAI22_X1 port map( A1 => n77_port, A2 => n11654, B1 => n205_port, 
                           B2 => n11637, ZN => n9417);
   U15289 : AOI21_X1 port map( B1 => n9432, B2 => n9433, A => n10841, ZN => 
                           n9431);
   U15290 : AOI221_X1 port map( B1 => n10795, B2 => n10391, C1 => n10778, C2 =>
                           n9943, A => n9435, ZN => n9432);
   U15291 : AOI221_X1 port map( B1 => n10830, B2 => n10392, C1 => n10812, C2 =>
                           n9944, A => n9434, ZN => n9433);
   U15292 : OAI22_X1 port map( A1 => n76_port, A2 => n11653, B1 => n204_port, 
                           B2 => n11636, ZN => n9435);
   U15293 : AOI21_X1 port map( B1 => n9450, B2 => n9451, A => n10841, ZN => 
                           n9449);
   U15294 : AOI221_X1 port map( B1 => n10795, B2 => n10393, C1 => n10778, C2 =>
                           n9945, A => n9453, ZN => n9450);
   U15295 : AOI221_X1 port map( B1 => n10830, B2 => n10394, C1 => n10812, C2 =>
                           n9946, A => n9452, ZN => n9451);
   U15296 : OAI22_X1 port map( A1 => n75_port, A2 => n11653, B1 => n203_port, 
                           B2 => n11636, ZN => n9453);
   U15297 : AOI21_X1 port map( B1 => n9468, B2 => n9469, A => n10841, ZN => 
                           n9467);
   U15298 : AOI221_X1 port map( B1 => n10795, B2 => n10395, C1 => n10778, C2 =>
                           n9947, A => n9471, ZN => n9468);
   U15299 : AOI221_X1 port map( B1 => n10831, B2 => n10396, C1 => n10813, C2 =>
                           n9948, A => n9470, ZN => n9469);
   U15300 : OAI22_X1 port map( A1 => n74_port, A2 => n11653, B1 => n202_port, 
                           B2 => n11636, ZN => n9471);
   U15301 : AOI21_X1 port map( B1 => n9486, B2 => n9487, A => n10841, ZN => 
                           n9485);
   U15302 : AOI221_X1 port map( B1 => n10795, B2 => n10397, C1 => n10778, C2 =>
                           n9949, A => n9489, ZN => n9486);
   U15303 : AOI221_X1 port map( B1 => n10831, B2 => n10398, C1 => n10813, C2 =>
                           n9950, A => n9488, ZN => n9487);
   U15304 : OAI22_X1 port map( A1 => n73_port, A2 => n11653, B1 => n201_port, 
                           B2 => n11636, ZN => n9489);
   U15305 : AOI21_X1 port map( B1 => n9504, B2 => n9505, A => n10841, ZN => 
                           n9503);
   U15306 : AOI221_X1 port map( B1 => n10795, B2 => n10399, C1 => n10778, C2 =>
                           n9951, A => n9507, ZN => n9504);
   U15307 : AOI221_X1 port map( B1 => n10831, B2 => n10400, C1 => n10813, C2 =>
                           n9952, A => n9506, ZN => n9505);
   U15308 : OAI22_X1 port map( A1 => n72_port, A2 => n11653, B1 => n200_port, 
                           B2 => n11636, ZN => n9507);
   U15309 : AOI21_X1 port map( B1 => n9522, B2 => n9523, A => n10841, ZN => 
                           n9521);
   U15310 : AOI221_X1 port map( B1 => n10795, B2 => n10401, C1 => n10778, C2 =>
                           n9953, A => n9525, ZN => n9522);
   U15311 : AOI221_X1 port map( B1 => n10831, B2 => n10402, C1 => n10813, C2 =>
                           n9954, A => n9524, ZN => n9523);
   U15312 : OAI22_X1 port map( A1 => n71_port, A2 => n11653, B1 => n199_port, 
                           B2 => n11636, ZN => n9525);
   U15313 : AOI21_X1 port map( B1 => n9540, B2 => n9541, A => n10841, ZN => 
                           n9539);
   U15314 : AOI221_X1 port map( B1 => n10796, B2 => n10403, C1 => n10779, C2 =>
                           n9955, A => n9543, ZN => n9540);
   U15315 : AOI221_X1 port map( B1 => n10831, B2 => n10404, C1 => n10813, C2 =>
                           n9956, A => n9542, ZN => n9541);
   U15316 : OAI22_X1 port map( A1 => n70_port, A2 => n11652, B1 => n198_port, 
                           B2 => n11635, ZN => n9543);
   U15317 : AOI21_X1 port map( B1 => n9558, B2 => n9559, A => n10841, ZN => 
                           n9557);
   U15318 : AOI221_X1 port map( B1 => n10796, B2 => n10405, C1 => n10779, C2 =>
                           n9957, A => n9561, ZN => n9558);
   U15319 : AOI221_X1 port map( B1 => n10831, B2 => n10406, C1 => n10813, C2 =>
                           n9958, A => n9560, ZN => n9559);
   U15320 : OAI22_X1 port map( A1 => n69_port, A2 => n11652, B1 => n197_port, 
                           B2 => n11635, ZN => n9561);
   U15321 : AOI21_X1 port map( B1 => n9576, B2 => n9577, A => n10841, ZN => 
                           n9575);
   U15322 : AOI221_X1 port map( B1 => n10796, B2 => n10407, C1 => n10779, C2 =>
                           n9959, A => n9579, ZN => n9576);
   U15323 : AOI221_X1 port map( B1 => n10832, B2 => n10408, C1 => n10814, C2 =>
                           n9960, A => n9578, ZN => n9577);
   U15324 : OAI22_X1 port map( A1 => n68_port, A2 => n11652, B1 => n196_port, 
                           B2 => n11635, ZN => n9579);
   U15325 : AOI21_X1 port map( B1 => n9594, B2 => n9595, A => n10841, ZN => 
                           n9593);
   U15326 : AOI221_X1 port map( B1 => n10796, B2 => n10409, C1 => n10779, C2 =>
                           n9961, A => n9597, ZN => n9594);
   U15327 : AOI221_X1 port map( B1 => n10832, B2 => n10410, C1 => n10814, C2 =>
                           n9962, A => n9596, ZN => n9595);
   U15328 : OAI22_X1 port map( A1 => n67_port, A2 => n11652, B1 => n195_port, 
                           B2 => n11635, ZN => n9597);
   U15329 : AOI21_X1 port map( B1 => n9612, B2 => n9613, A => n10841, ZN => 
                           n9611);
   U15330 : AOI221_X1 port map( B1 => n10796, B2 => n10411, C1 => n10779, C2 =>
                           n9963, A => n9615, ZN => n9612);
   U15331 : AOI221_X1 port map( B1 => n10832, B2 => n10412, C1 => n10814, C2 =>
                           n9964, A => n9614, ZN => n9613);
   U15332 : OAI22_X1 port map( A1 => n66_port, A2 => n11652, B1 => n194_port, 
                           B2 => n11635, ZN => n9615);
   U15333 : AOI21_X1 port map( B1 => n9630, B2 => n9631, A => n10841, ZN => 
                           n9629);
   U15334 : AOI221_X1 port map( B1 => n10796, B2 => n10413, C1 => n10779, C2 =>
                           n9965, A => n9633, ZN => n9630);
   U15335 : AOI221_X1 port map( B1 => n10832, B2 => n10414, C1 => n10814, C2 =>
                           n9966, A => n9632, ZN => n9631);
   U15336 : OAI22_X1 port map( A1 => n65_port, A2 => n11652, B1 => n193_port, 
                           B2 => n11635, ZN => n9633);
   U15337 : AOI21_X1 port map( B1 => n7303, B2 => n7304, A => n10992, ZN => 
                           n7292);
   U15338 : AOI221_X1 port map( B1 => n11012, B2 => n10415, C1 => n10995, C2 =>
                           n9967, A => n7307, ZN => n7303);
   U15339 : AOI221_X1 port map( B1 => n11047, B2 => n10416, C1 => n11029, C2 =>
                           n9968, A => n7306, ZN => n7304);
   U15340 : OAI22_X1 port map( A1 => n640_port, A2 => n11594, B1 => n768_port, 
                           B2 => n11577, ZN => n7307);
   U15341 : AOI21_X1 port map( B1 => n7338, B2 => n7339, A => n10992, ZN => 
                           n7332);
   U15342 : AOI221_X1 port map( B1 => n11012, B2 => n10417, C1 => n10995, C2 =>
                           n9969, A => n7341, ZN => n7338);
   U15343 : AOI221_X1 port map( B1 => n11047, B2 => n10418, C1 => n11029, C2 =>
                           n9970, A => n7340, ZN => n7339);
   U15344 : OAI22_X1 port map( A1 => n639_port, A2 => n11594, B1 => n767_port, 
                           B2 => n11577, ZN => n7341);
   U15345 : AOI21_X1 port map( B1 => n7356, B2 => n7357, A => n10992, ZN => 
                           n7350);
   U15346 : AOI221_X1 port map( B1 => n11012, B2 => n10419, C1 => n10995, C2 =>
                           n9971, A => n7359, ZN => n7356);
   U15347 : AOI221_X1 port map( B1 => n11047, B2 => n10420, C1 => n11029, C2 =>
                           n9972, A => n7358, ZN => n7357);
   U15348 : OAI22_X1 port map( A1 => n638_port, A2 => n11594, B1 => n766_port, 
                           B2 => n11577, ZN => n7359);
   U15349 : AOI21_X1 port map( B1 => n7374, B2 => n7375, A => n10992, ZN => 
                           n7368);
   U15350 : AOI221_X1 port map( B1 => n11012, B2 => n10421, C1 => n10995, C2 =>
                           n9973, A => n7377, ZN => n7374);
   U15351 : AOI221_X1 port map( B1 => n11047, B2 => n10422, C1 => n11029, C2 =>
                           n9974, A => n7376, ZN => n7375);
   U15352 : OAI22_X1 port map( A1 => n637_port, A2 => n11594, B1 => n765_port, 
                           B2 => n11577, ZN => n7377);
   U15353 : AOI21_X1 port map( B1 => n7392, B2 => n7393, A => n10991, ZN => 
                           n7386);
   U15354 : AOI221_X1 port map( B1 => n11012, B2 => n10423, C1 => n10995, C2 =>
                           n9975, A => n7395, ZN => n7392);
   U15355 : AOI221_X1 port map( B1 => n11047, B2 => n10424, C1 => n11029, C2 =>
                           n9976, A => n7394, ZN => n7393);
   U15356 : OAI22_X1 port map( A1 => n636_port, A2 => n11593, B1 => n764_port, 
                           B2 => n11576, ZN => n7395);
   U15357 : AOI21_X1 port map( B1 => n7410, B2 => n7411, A => n10991, ZN => 
                           n7404);
   U15358 : AOI221_X1 port map( B1 => n11012, B2 => n10425, C1 => n10995, C2 =>
                           n9977, A => n7413, ZN => n7410);
   U15359 : AOI221_X1 port map( B1 => n11047, B2 => n10426, C1 => n11029, C2 =>
                           n9978, A => n7412, ZN => n7411);
   U15360 : OAI22_X1 port map( A1 => n635_port, A2 => n11593, B1 => n763_port, 
                           B2 => n11576, ZN => n7413);
   U15361 : AOI21_X1 port map( B1 => n7428, B2 => n7429, A => n10991, ZN => 
                           n7422);
   U15362 : AOI221_X1 port map( B1 => n11013, B2 => n10427, C1 => n10996, C2 =>
                           n9979, A => n7431, ZN => n7428);
   U15363 : AOI221_X1 port map( B1 => n11048, B2 => n10428, C1 => n11030, C2 =>
                           n9980, A => n7430, ZN => n7429);
   U15364 : OAI22_X1 port map( A1 => n634_port, A2 => n11593, B1 => n762_port, 
                           B2 => n11576, ZN => n7431);
   U15365 : AOI21_X1 port map( B1 => n7446, B2 => n7447, A => n10991, ZN => 
                           n7440);
   U15366 : AOI221_X1 port map( B1 => n11013, B2 => n10429, C1 => n10996, C2 =>
                           n9981, A => n7449, ZN => n7446);
   U15367 : AOI221_X1 port map( B1 => n11048, B2 => n10430, C1 => n11030, C2 =>
                           n9982, A => n7448, ZN => n7447);
   U15368 : OAI22_X1 port map( A1 => n633_port, A2 => n11593, B1 => n761_port, 
                           B2 => n11576, ZN => n7449);
   U15369 : AOI21_X1 port map( B1 => n7464, B2 => n7465, A => n10991, ZN => 
                           n7458);
   U15370 : AOI221_X1 port map( B1 => n11013, B2 => n10431, C1 => n10996, C2 =>
                           n9983, A => n7467, ZN => n7464);
   U15371 : AOI221_X1 port map( B1 => n11048, B2 => n10432, C1 => n11030, C2 =>
                           n9984, A => n7466, ZN => n7465);
   U15372 : OAI22_X1 port map( A1 => n632_port, A2 => n11593, B1 => n760_port, 
                           B2 => n11576, ZN => n7467);
   U15373 : AOI21_X1 port map( B1 => n7482, B2 => n7483, A => n10991, ZN => 
                           n7476);
   U15374 : AOI221_X1 port map( B1 => n11013, B2 => n10433, C1 => n10996, C2 =>
                           n9985, A => n7485, ZN => n7482);
   U15375 : AOI221_X1 port map( B1 => n11048, B2 => n10434, C1 => n11030, C2 =>
                           n9986, A => n7484, ZN => n7483);
   U15376 : OAI22_X1 port map( A1 => n631_port, A2 => n11593, B1 => n759_port, 
                           B2 => n11576, ZN => n7485);
   U15377 : AOI21_X1 port map( B1 => n7500, B2 => n7501, A => n10991, ZN => 
                           n7494);
   U15378 : AOI221_X1 port map( B1 => n11013, B2 => n10435, C1 => n10996, C2 =>
                           n9987, A => n7503, ZN => n7500);
   U15379 : AOI221_X1 port map( B1 => n11048, B2 => n10436, C1 => n11030, C2 =>
                           n9988, A => n7502, ZN => n7501);
   U15380 : OAI22_X1 port map( A1 => n630_port, A2 => n11592, B1 => n758_port, 
                           B2 => n11575, ZN => n7503);
   U15381 : AOI21_X1 port map( B1 => n7518, B2 => n7519, A => n10991, ZN => 
                           n7512);
   U15382 : AOI221_X1 port map( B1 => n11013, B2 => n10437, C1 => n10996, C2 =>
                           n9989, A => n7521, ZN => n7518);
   U15383 : AOI221_X1 port map( B1 => n11048, B2 => n10438, C1 => n11030, C2 =>
                           n9990, A => n7520, ZN => n7519);
   U15384 : OAI22_X1 port map( A1 => n629_port, A2 => n11592, B1 => n757_port, 
                           B2 => n11575, ZN => n7521);
   U15385 : AOI21_X1 port map( B1 => n7536, B2 => n7537, A => n10991, ZN => 
                           n7530);
   U15386 : AOI221_X1 port map( B1 => n11013, B2 => n10439, C1 => n10996, C2 =>
                           n9991, A => n7539, ZN => n7536);
   U15387 : AOI221_X1 port map( B1 => n11049, B2 => n10440, C1 => n11031, C2 =>
                           n9992, A => n7538, ZN => n7537);
   U15388 : OAI22_X1 port map( A1 => n628_port, A2 => n11592, B1 => n756_port, 
                           B2 => n11575, ZN => n7539);
   U15389 : AOI21_X1 port map( B1 => n7554, B2 => n7555, A => n10991, ZN => 
                           n7548);
   U15390 : AOI221_X1 port map( B1 => n11014, B2 => n10441, C1 => n10997, C2 =>
                           n9993, A => n7557, ZN => n7554);
   U15391 : AOI221_X1 port map( B1 => n11049, B2 => n10442, C1 => n11031, C2 =>
                           n9994, A => n7556, ZN => n7555);
   U15392 : OAI22_X1 port map( A1 => n627_port, A2 => n11592, B1 => n755_port, 
                           B2 => n11575, ZN => n7557);
   U15393 : AOI21_X1 port map( B1 => n7572, B2 => n7573, A => n10991, ZN => 
                           n7566);
   U15394 : AOI221_X1 port map( B1 => n11014, B2 => n10443, C1 => n10997, C2 =>
                           n9995, A => n7575, ZN => n7572);
   U15395 : AOI221_X1 port map( B1 => n11049, B2 => n10444, C1 => n11031, C2 =>
                           n9996, A => n7574, ZN => n7573);
   U15396 : OAI22_X1 port map( A1 => n626_port, A2 => n11592, B1 => n754_port, 
                           B2 => n11575, ZN => n7575);
   U15397 : AOI21_X1 port map( B1 => n7590, B2 => n7591, A => n10991, ZN => 
                           n7584);
   U15398 : AOI221_X1 port map( B1 => n11014, B2 => n10445, C1 => n10997, C2 =>
                           n9997, A => n7593, ZN => n7590);
   U15399 : AOI221_X1 port map( B1 => n11049, B2 => n10446, C1 => n11031, C2 =>
                           n9998, A => n7592, ZN => n7591);
   U15400 : OAI22_X1 port map( A1 => n625_port, A2 => n11592, B1 => n753_port, 
                           B2 => n11575, ZN => n7593);
   U15401 : AOI21_X1 port map( B1 => n7608, B2 => n7609, A => n10990, ZN => 
                           n7602);
   U15402 : AOI221_X1 port map( B1 => n11014, B2 => n10447, C1 => n10997, C2 =>
                           n9999, A => n7611, ZN => n7608);
   U15403 : AOI221_X1 port map( B1 => n11049, B2 => n10448, C1 => n11031, C2 =>
                           n10000, A => n7610, ZN => n7609);
   U15404 : OAI22_X1 port map( A1 => n624_port, A2 => n11591, B1 => n752_port, 
                           B2 => n11574, ZN => n7611);
   U15405 : AOI21_X1 port map( B1 => n7626, B2 => n7627, A => n10990, ZN => 
                           n7620);
   U15406 : AOI221_X1 port map( B1 => n11014, B2 => n10449, C1 => n10997, C2 =>
                           n10001, A => n7629, ZN => n7626);
   U15407 : AOI221_X1 port map( B1 => n11049, B2 => n10450, C1 => n11031, C2 =>
                           n10002, A => n7628, ZN => n7627);
   U15408 : OAI22_X1 port map( A1 => n623_port, A2 => n11591, B1 => n751_port, 
                           B2 => n11574, ZN => n7629);
   U15409 : AOI21_X1 port map( B1 => n7644, B2 => n7645, A => n10990, ZN => 
                           n7638);
   U15410 : AOI221_X1 port map( B1 => n11014, B2 => n10451, C1 => n10997, C2 =>
                           n10003, A => n7647, ZN => n7644);
   U15411 : AOI221_X1 port map( B1 => n11050, B2 => n10452, C1 => n11032, C2 =>
                           n10004, A => n7646, ZN => n7645);
   U15412 : OAI22_X1 port map( A1 => n622_port, A2 => n11591, B1 => n750_port, 
                           B2 => n11574, ZN => n7647);
   U15413 : AOI21_X1 port map( B1 => n7662, B2 => n7663, A => n10990, ZN => 
                           n7656);
   U15414 : AOI221_X1 port map( B1 => n11015, B2 => n10453, C1 => n10998, C2 =>
                           n10005, A => n7665, ZN => n7662);
   U15415 : AOI221_X1 port map( B1 => n11050, B2 => n10454, C1 => n11032, C2 =>
                           n10006, A => n7664, ZN => n7663);
   U15416 : OAI22_X1 port map( A1 => n621_port, A2 => n11591, B1 => n749_port, 
                           B2 => n11574, ZN => n7665);
   U15417 : AOI21_X1 port map( B1 => n7680, B2 => n7681, A => n10990, ZN => 
                           n7674);
   U15418 : AOI221_X1 port map( B1 => n11015, B2 => n10455, C1 => n10998, C2 =>
                           n10007, A => n7683, ZN => n7680);
   U15419 : AOI221_X1 port map( B1 => n11050, B2 => n10456, C1 => n11032, C2 =>
                           n10008, A => n7682, ZN => n7681);
   U15420 : OAI22_X1 port map( A1 => n620_port, A2 => n11591, B1 => n748_port, 
                           B2 => n11574, ZN => n7683);
   U15421 : AOI21_X1 port map( B1 => n7698, B2 => n7699, A => n10990, ZN => 
                           n7692);
   U15422 : AOI221_X1 port map( B1 => n11015, B2 => n10457, C1 => n10998, C2 =>
                           n10009, A => n7701, ZN => n7698);
   U15423 : AOI221_X1 port map( B1 => n11050, B2 => n10458, C1 => n11032, C2 =>
                           n10010, A => n7700, ZN => n7699);
   U15424 : OAI22_X1 port map( A1 => n619_port, A2 => n11591, B1 => n747_port, 
                           B2 => n11574, ZN => n7701);
   U15425 : AOI21_X1 port map( B1 => n7716, B2 => n7717, A => n10990, ZN => 
                           n7710);
   U15426 : AOI221_X1 port map( B1 => n11015, B2 => n10459, C1 => n10998, C2 =>
                           n10011, A => n7719, ZN => n7716);
   U15427 : AOI221_X1 port map( B1 => n11050, B2 => n10460, C1 => n11032, C2 =>
                           n10012, A => n7718, ZN => n7717);
   U15428 : OAI22_X1 port map( A1 => n618_port, A2 => n11590, B1 => n746_port, 
                           B2 => n11573, ZN => n7719);
   U15429 : AOI21_X1 port map( B1 => n7734, B2 => n7735, A => n10990, ZN => 
                           n7728);
   U15430 : AOI221_X1 port map( B1 => n11015, B2 => n10461, C1 => n10998, C2 =>
                           n10013, A => n7737, ZN => n7734);
   U15431 : AOI221_X1 port map( B1 => n11050, B2 => n10462, C1 => n11032, C2 =>
                           n10014, A => n7736, ZN => n7735);
   U15432 : OAI22_X1 port map( A1 => n617_port, A2 => n11590, B1 => n745_port, 
                           B2 => n11573, ZN => n7737);
   U15433 : AOI21_X1 port map( B1 => n7752, B2 => n7753, A => n10990, ZN => 
                           n7746);
   U15434 : AOI221_X1 port map( B1 => n11015, B2 => n10463, C1 => n10998, C2 =>
                           n10015, A => n7755, ZN => n7752);
   U15435 : AOI221_X1 port map( B1 => n11051, B2 => n10464, C1 => n11033, C2 =>
                           n10016, A => n7754, ZN => n7753);
   U15436 : OAI22_X1 port map( A1 => n616_port, A2 => n11590, B1 => n744_port, 
                           B2 => n11573, ZN => n7755);
   U15437 : AOI21_X1 port map( B1 => n7770, B2 => n7771, A => n10990, ZN => 
                           n7764);
   U15438 : AOI221_X1 port map( B1 => n11015, B2 => n10465, C1 => n10998, C2 =>
                           n10017, A => n7773, ZN => n7770);
   U15439 : AOI221_X1 port map( B1 => n11051, B2 => n10466, C1 => n11033, C2 =>
                           n10018, A => n7772, ZN => n7771);
   U15440 : OAI22_X1 port map( A1 => n615_port, A2 => n11590, B1 => n743_port, 
                           B2 => n11573, ZN => n7773);
   U15441 : AOI21_X1 port map( B1 => n7788, B2 => n7789, A => n10990, ZN => 
                           n7782);
   U15442 : AOI221_X1 port map( B1 => n11016, B2 => n10467, C1 => n10999, C2 =>
                           n10019, A => n7791, ZN => n7788);
   U15443 : AOI221_X1 port map( B1 => n11051, B2 => n10468, C1 => n11033, C2 =>
                           n10020, A => n7790, ZN => n7789);
   U15444 : OAI22_X1 port map( A1 => n614_port, A2 => n11590, B1 => n742_port, 
                           B2 => n11573, ZN => n7791);
   U15445 : AOI21_X1 port map( B1 => n7806, B2 => n7807, A => n10990, ZN => 
                           n7800);
   U15446 : AOI221_X1 port map( B1 => n11016, B2 => n10469, C1 => n10999, C2 =>
                           n10021, A => n7809, ZN => n7806);
   U15447 : AOI221_X1 port map( B1 => n11051, B2 => n10470, C1 => n11033, C2 =>
                           n10022, A => n7808, ZN => n7807);
   U15448 : OAI22_X1 port map( A1 => n613_port, A2 => n11590, B1 => n741_port, 
                           B2 => n11573, ZN => n7809);
   U15449 : AOI21_X1 port map( B1 => n7824, B2 => n7825, A => n10989, ZN => 
                           n7818);
   U15450 : AOI221_X1 port map( B1 => n11016, B2 => n10471, C1 => n10999, C2 =>
                           n10023, A => n7827, ZN => n7824);
   U15451 : AOI221_X1 port map( B1 => n11051, B2 => n10472, C1 => n11033, C2 =>
                           n10024, A => n7826, ZN => n7825);
   U15452 : OAI22_X1 port map( A1 => n612_port, A2 => n11589, B1 => n740_port, 
                           B2 => n11572, ZN => n7827);
   U15453 : AOI21_X1 port map( B1 => n7842, B2 => n7843, A => n10989, ZN => 
                           n7836);
   U15454 : AOI221_X1 port map( B1 => n11016, B2 => n10473, C1 => n10999, C2 =>
                           n10025, A => n7845, ZN => n7842);
   U15455 : AOI221_X1 port map( B1 => n11051, B2 => n10474, C1 => n11033, C2 =>
                           n10026, A => n7844, ZN => n7843);
   U15456 : OAI22_X1 port map( A1 => n611_port, A2 => n11589, B1 => n739_port, 
                           B2 => n11572, ZN => n7845);
   U15457 : AOI21_X1 port map( B1 => n7860, B2 => n7861, A => n10989, ZN => 
                           n7854);
   U15458 : AOI221_X1 port map( B1 => n11016, B2 => n10475, C1 => n10999, C2 =>
                           n10027, A => n7863, ZN => n7860);
   U15459 : AOI221_X1 port map( B1 => n11052, B2 => n10476, C1 => n11034, C2 =>
                           n10028, A => n7862, ZN => n7861);
   U15460 : OAI22_X1 port map( A1 => n610_port, A2 => n11589, B1 => n738_port, 
                           B2 => n11572, ZN => n7863);
   U15461 : AOI21_X1 port map( B1 => n7878, B2 => n7879, A => n10989, ZN => 
                           n7872);
   U15462 : AOI221_X1 port map( B1 => n11016, B2 => n10477, C1 => n10999, C2 =>
                           n10029, A => n7881, ZN => n7878);
   U15463 : AOI221_X1 port map( B1 => n11052, B2 => n10478, C1 => n11034, C2 =>
                           n10030, A => n7880, ZN => n7879);
   U15464 : OAI22_X1 port map( A1 => n609_port, A2 => n11589, B1 => n737_port, 
                           B2 => n11572, ZN => n7881);
   U15465 : AOI21_X1 port map( B1 => n7896, B2 => n7897, A => n10989, ZN => 
                           n7890);
   U15466 : AOI221_X1 port map( B1 => n11017, B2 => n10479, C1 => n11000, C2 =>
                           n10031, A => n7899, ZN => n7896);
   U15467 : AOI221_X1 port map( B1 => n11052, B2 => n10480, C1 => n11034, C2 =>
                           n10032, A => n7898, ZN => n7897);
   U15468 : OAI22_X1 port map( A1 => n608_port, A2 => n11589, B1 => n736_port, 
                           B2 => n11572, ZN => n7899);
   U15469 : AOI21_X1 port map( B1 => n7914, B2 => n7915, A => n10989, ZN => 
                           n7908);
   U15470 : AOI221_X1 port map( B1 => n11017, B2 => n10481, C1 => n11000, C2 =>
                           n10033, A => n7917, ZN => n7914);
   U15471 : AOI221_X1 port map( B1 => n11052, B2 => n10482, C1 => n11034, C2 =>
                           n10034, A => n7916, ZN => n7915);
   U15472 : OAI22_X1 port map( A1 => n607_port, A2 => n11589, B1 => n735_port, 
                           B2 => n11572, ZN => n7917);
   U15473 : AOI21_X1 port map( B1 => n7932, B2 => n7933, A => n10989, ZN => 
                           n7926);
   U15474 : AOI221_X1 port map( B1 => n11017, B2 => n10483, C1 => n11000, C2 =>
                           n10035, A => n7935, ZN => n7932);
   U15475 : AOI221_X1 port map( B1 => n11052, B2 => n10484, C1 => n11034, C2 =>
                           n10036, A => n7934, ZN => n7933);
   U15476 : OAI22_X1 port map( A1 => n606_port, A2 => n11588, B1 => n734_port, 
                           B2 => n11571, ZN => n7935);
   U15477 : AOI21_X1 port map( B1 => n7950, B2 => n7951, A => n10989, ZN => 
                           n7944);
   U15478 : AOI221_X1 port map( B1 => n11017, B2 => n10485, C1 => n11000, C2 =>
                           n10037, A => n7953, ZN => n7950);
   U15479 : AOI221_X1 port map( B1 => n11052, B2 => n10486, C1 => n11034, C2 =>
                           n10038, A => n7952, ZN => n7951);
   U15480 : OAI22_X1 port map( A1 => n605_port, A2 => n11588, B1 => n733_port, 
                           B2 => n11571, ZN => n7953);
   U15481 : AOI21_X1 port map( B1 => n7968, B2 => n7969, A => n10989, ZN => 
                           n7962);
   U15482 : AOI221_X1 port map( B1 => n11017, B2 => n10487, C1 => n11000, C2 =>
                           n10039, A => n7971, ZN => n7968);
   U15483 : AOI221_X1 port map( B1 => n11053, B2 => n10488, C1 => n11035, C2 =>
                           n10040, A => n7970, ZN => n7969);
   U15484 : OAI22_X1 port map( A1 => n604_port, A2 => n11588, B1 => n732_port, 
                           B2 => n11571, ZN => n7971);
   U15485 : AOI21_X1 port map( B1 => n7986, B2 => n7987, A => n10989, ZN => 
                           n7980);
   U15486 : AOI221_X1 port map( B1 => n11017, B2 => n10489, C1 => n11000, C2 =>
                           n10041, A => n7989, ZN => n7986);
   U15487 : AOI221_X1 port map( B1 => n11053, B2 => n10490, C1 => n11035, C2 =>
                           n10042, A => n7988, ZN => n7987);
   U15488 : OAI22_X1 port map( A1 => n603_port, A2 => n11588, B1 => n731_port, 
                           B2 => n11571, ZN => n7989);
   U15489 : AOI21_X1 port map( B1 => n8004, B2 => n8005, A => n10989, ZN => 
                           n7998);
   U15490 : AOI221_X1 port map( B1 => n11018, B2 => n10491, C1 => n11001, C2 =>
                           n10043, A => n8007, ZN => n8004);
   U15491 : AOI221_X1 port map( B1 => n11053, B2 => n10492, C1 => n11035, C2 =>
                           n10044, A => n8006, ZN => n8005);
   U15492 : OAI22_X1 port map( A1 => n602_port, A2 => n11588, B1 => n730_port, 
                           B2 => n11571, ZN => n8007);
   U15493 : AOI21_X1 port map( B1 => n8022, B2 => n8023, A => n10989, ZN => 
                           n8016);
   U15494 : AOI221_X1 port map( B1 => n11018, B2 => n10493, C1 => n11001, C2 =>
                           n10045, A => n8025, ZN => n8022);
   U15495 : AOI221_X1 port map( B1 => n11053, B2 => n10494, C1 => n11035, C2 =>
                           n10046, A => n8024, ZN => n8023);
   U15496 : OAI22_X1 port map( A1 => n601_port, A2 => n11588, B1 => n729_port, 
                           B2 => n11571, ZN => n8025);
   U15497 : AOI21_X1 port map( B1 => n8040, B2 => n8041, A => n10988, ZN => 
                           n8034);
   U15498 : AOI221_X1 port map( B1 => n11018, B2 => n10495, C1 => n11001, C2 =>
                           n10047, A => n8043, ZN => n8040);
   U15499 : AOI221_X1 port map( B1 => n11053, B2 => n10496, C1 => n11035, C2 =>
                           n10048, A => n8042, ZN => n8041);
   U15500 : OAI22_X1 port map( A1 => n600_port, A2 => n11587, B1 => n728_port, 
                           B2 => n11570, ZN => n8043);
   U15501 : AOI21_X1 port map( B1 => n8058, B2 => n8059, A => n10988, ZN => 
                           n8052);
   U15502 : AOI221_X1 port map( B1 => n11018, B2 => n10497, C1 => n11001, C2 =>
                           n10049, A => n8061, ZN => n8058);
   U15503 : AOI221_X1 port map( B1 => n11053, B2 => n10498, C1 => n11035, C2 =>
                           n10050, A => n8060, ZN => n8059);
   U15504 : OAI22_X1 port map( A1 => n599_port, A2 => n11587, B1 => n727_port, 
                           B2 => n11570, ZN => n8061);
   U15505 : AOI21_X1 port map( B1 => n8076, B2 => n8077, A => n10988, ZN => 
                           n8070);
   U15506 : AOI221_X1 port map( B1 => n11018, B2 => n10499, C1 => n11001, C2 =>
                           n10051, A => n8079, ZN => n8076);
   U15507 : AOI221_X1 port map( B1 => n11054, B2 => n10500, C1 => n11036, C2 =>
                           n10052, A => n8078, ZN => n8077);
   U15508 : OAI22_X1 port map( A1 => n598_port, A2 => n11587, B1 => n726_port, 
                           B2 => n11570, ZN => n8079);
   U15509 : AOI21_X1 port map( B1 => n8094, B2 => n8095, A => n10988, ZN => 
                           n8088);
   U15510 : AOI221_X1 port map( B1 => n11018, B2 => n10501, C1 => n11001, C2 =>
                           n10053, A => n8097, ZN => n8094);
   U15511 : AOI221_X1 port map( B1 => n11054, B2 => n10502, C1 => n11036, C2 =>
                           n10054, A => n8096, ZN => n8095);
   U15512 : OAI22_X1 port map( A1 => n597_port, A2 => n11587, B1 => n725_port, 
                           B2 => n11570, ZN => n8097);
   U15513 : AOI21_X1 port map( B1 => n8112, B2 => n8113, A => n10988, ZN => 
                           n8106);
   U15514 : AOI221_X1 port map( B1 => n11018, B2 => n10503, C1 => n11001, C2 =>
                           n10055, A => n8115, ZN => n8112);
   U15515 : AOI221_X1 port map( B1 => n11054, B2 => n10504, C1 => n11036, C2 =>
                           n10056, A => n8114, ZN => n8113);
   U15516 : OAI22_X1 port map( A1 => n596_port, A2 => n11587, B1 => n724_port, 
                           B2 => n11570, ZN => n8115);
   U15517 : AOI21_X1 port map( B1 => n8130, B2 => n8131, A => n10988, ZN => 
                           n8124);
   U15518 : AOI221_X1 port map( B1 => n11019, B2 => n10505, C1 => n11002, C2 =>
                           n10057, A => n8133, ZN => n8130);
   U15519 : AOI221_X1 port map( B1 => n11054, B2 => n10506, C1 => n11036, C2 =>
                           n10058, A => n8132, ZN => n8131);
   U15520 : OAI22_X1 port map( A1 => n595_port, A2 => n11587, B1 => n723_port, 
                           B2 => n11570, ZN => n8133);
   U15521 : AOI21_X1 port map( B1 => n8148, B2 => n8149, A => n10988, ZN => 
                           n8142);
   U15522 : AOI221_X1 port map( B1 => n11019, B2 => n10507, C1 => n11002, C2 =>
                           n10059, A => n8151, ZN => n8148);
   U15523 : AOI221_X1 port map( B1 => n11054, B2 => n10508, C1 => n11036, C2 =>
                           n10060, A => n8150, ZN => n8149);
   U15524 : OAI22_X1 port map( A1 => n594_port, A2 => n11586, B1 => n722_port, 
                           B2 => n11569, ZN => n8151);
   U15525 : AOI21_X1 port map( B1 => n8166, B2 => n8167, A => n10988, ZN => 
                           n8160);
   U15526 : AOI221_X1 port map( B1 => n11019, B2 => n10509, C1 => n11002, C2 =>
                           n10061, A => n8169, ZN => n8166);
   U15527 : AOI221_X1 port map( B1 => n11054, B2 => n10510, C1 => n11036, C2 =>
                           n10062, A => n8168, ZN => n8167);
   U15528 : OAI22_X1 port map( A1 => n593_port, A2 => n11586, B1 => n721_port, 
                           B2 => n11569, ZN => n8169);
   U15529 : AOI21_X1 port map( B1 => n8184, B2 => n8185, A => n10988, ZN => 
                           n8178);
   U15530 : AOI221_X1 port map( B1 => n11019, B2 => n10511, C1 => n11002, C2 =>
                           n10063, A => n8187, ZN => n8184);
   U15531 : AOI221_X1 port map( B1 => n11055, B2 => n10512, C1 => n11037, C2 =>
                           n10064, A => n8186, ZN => n8185);
   U15532 : OAI22_X1 port map( A1 => n592_port, A2 => n11586, B1 => n720_port, 
                           B2 => n11569, ZN => n8187);
   U15533 : AOI21_X1 port map( B1 => n8202, B2 => n8203, A => n10988, ZN => 
                           n8196);
   U15534 : AOI221_X1 port map( B1 => n11019, B2 => n10513, C1 => n11002, C2 =>
                           n10065, A => n8205, ZN => n8202);
   U15535 : AOI221_X1 port map( B1 => n11055, B2 => n10514, C1 => n11037, C2 =>
                           n10066, A => n8204, ZN => n8203);
   U15536 : OAI22_X1 port map( A1 => n591_port, A2 => n11586, B1 => n719_port, 
                           B2 => n11569, ZN => n8205);
   U15537 : AOI21_X1 port map( B1 => n8220, B2 => n8221, A => n10988, ZN => 
                           n8214);
   U15538 : AOI221_X1 port map( B1 => n11019, B2 => n10515, C1 => n11002, C2 =>
                           n10067, A => n8223, ZN => n8220);
   U15539 : AOI221_X1 port map( B1 => n11055, B2 => n10516, C1 => n11037, C2 =>
                           n10068, A => n8222, ZN => n8221);
   U15540 : OAI22_X1 port map( A1 => n590_port, A2 => n11586, B1 => n718_port, 
                           B2 => n11569, ZN => n8223);
   U15541 : AOI21_X1 port map( B1 => n8238, B2 => n8239, A => n10988, ZN => 
                           n8232);
   U15542 : AOI221_X1 port map( B1 => n11020, B2 => n10517, C1 => n11003, C2 =>
                           n10069, A => n8241, ZN => n8238);
   U15543 : AOI221_X1 port map( B1 => n11055, B2 => n10518, C1 => n11037, C2 =>
                           n10070, A => n8240, ZN => n8239);
   U15544 : OAI22_X1 port map( A1 => n589_port, A2 => n11586, B1 => n717_port, 
                           B2 => n11569, ZN => n8241);
   U15545 : AOI21_X1 port map( B1 => n8256, B2 => n8257, A => n10987, ZN => 
                           n8250);
   U15546 : AOI221_X1 port map( B1 => n11020, B2 => n10519, C1 => n11003, C2 =>
                           n10071, A => n8259, ZN => n8256);
   U15547 : AOI221_X1 port map( B1 => n11055, B2 => n10520, C1 => n11037, C2 =>
                           n10072, A => n8258, ZN => n8257);
   U15548 : OAI22_X1 port map( A1 => n588_port, A2 => n11585, B1 => n716_port, 
                           B2 => n11568, ZN => n8259);
   U15549 : AOI21_X1 port map( B1 => n8274, B2 => n8275, A => n10987, ZN => 
                           n8268);
   U15550 : AOI221_X1 port map( B1 => n11020, B2 => n10521, C1 => n11003, C2 =>
                           n10073, A => n8277, ZN => n8274);
   U15551 : AOI221_X1 port map( B1 => n11055, B2 => n10522, C1 => n11037, C2 =>
                           n10074, A => n8276, ZN => n8275);
   U15552 : OAI22_X1 port map( A1 => n587_port, A2 => n11585, B1 => n715_port, 
                           B2 => n11568, ZN => n8277);
   U15553 : AOI21_X1 port map( B1 => n8292, B2 => n8293, A => n10987, ZN => 
                           n8286);
   U15554 : AOI221_X1 port map( B1 => n11020, B2 => n10523, C1 => n11003, C2 =>
                           n10075, A => n8295, ZN => n8292);
   U15555 : AOI221_X1 port map( B1 => n11056, B2 => n10524, C1 => n11038, C2 =>
                           n10076, A => n8294, ZN => n8293);
   U15556 : OAI22_X1 port map( A1 => n586_port, A2 => n11585, B1 => n714_port, 
                           B2 => n11568, ZN => n8295);
   U15557 : AOI21_X1 port map( B1 => n8310, B2 => n8311, A => n10987, ZN => 
                           n8304);
   U15558 : AOI221_X1 port map( B1 => n11020, B2 => n10525, C1 => n11003, C2 =>
                           n10077, A => n8313, ZN => n8310);
   U15559 : AOI221_X1 port map( B1 => n11056, B2 => n10526, C1 => n11038, C2 =>
                           n10078, A => n8312, ZN => n8311);
   U15560 : OAI22_X1 port map( A1 => n585_port, A2 => n11585, B1 => n713_port, 
                           B2 => n11568, ZN => n8313);
   U15561 : AOI21_X1 port map( B1 => n8328, B2 => n8329, A => n10987, ZN => 
                           n8322);
   U15562 : AOI221_X1 port map( B1 => n11020, B2 => n10527, C1 => n11003, C2 =>
                           n10079, A => n8331, ZN => n8328);
   U15563 : AOI221_X1 port map( B1 => n11056, B2 => n10528, C1 => n11038, C2 =>
                           n10080, A => n8330, ZN => n8329);
   U15564 : OAI22_X1 port map( A1 => n584_port, A2 => n11585, B1 => n712_port, 
                           B2 => n11568, ZN => n8331);
   U15565 : AOI21_X1 port map( B1 => n8346, B2 => n8347, A => n10987, ZN => 
                           n8340);
   U15566 : AOI221_X1 port map( B1 => n11020, B2 => n10529, C1 => n11003, C2 =>
                           n10081, A => n8349, ZN => n8346);
   U15567 : AOI221_X1 port map( B1 => n11056, B2 => n10530, C1 => n11038, C2 =>
                           n10082, A => n8348, ZN => n8347);
   U15568 : OAI22_X1 port map( A1 => n583_port, A2 => n11585, B1 => n711_port, 
                           B2 => n11568, ZN => n8349);
   U15569 : AOI21_X1 port map( B1 => n8364, B2 => n8365, A => n10987, ZN => 
                           n8358);
   U15570 : AOI221_X1 port map( B1 => n11021, B2 => n10531, C1 => n11004, C2 =>
                           n10083, A => n8367, ZN => n8364);
   U15571 : AOI221_X1 port map( B1 => n11056, B2 => n10532, C1 => n11038, C2 =>
                           n10084, A => n8366, ZN => n8365);
   U15572 : OAI22_X1 port map( A1 => n582_port, A2 => n11584, B1 => n710_port, 
                           B2 => n11567, ZN => n8367);
   U15573 : AOI21_X1 port map( B1 => n8382, B2 => n8383, A => n10987, ZN => 
                           n8376);
   U15574 : AOI221_X1 port map( B1 => n11021, B2 => n10533, C1 => n11004, C2 =>
                           n10085, A => n8385, ZN => n8382);
   U15575 : AOI221_X1 port map( B1 => n11056, B2 => n10534, C1 => n11038, C2 =>
                           n10086, A => n8384, ZN => n8383);
   U15576 : OAI22_X1 port map( A1 => n581_port, A2 => n11584, B1 => n709_port, 
                           B2 => n11567, ZN => n8385);
   U15577 : AOI21_X1 port map( B1 => n8400, B2 => n8401, A => n10987, ZN => 
                           n8394);
   U15578 : AOI221_X1 port map( B1 => n11021, B2 => n10535, C1 => n11004, C2 =>
                           n10087, A => n8403, ZN => n8400);
   U15579 : AOI221_X1 port map( B1 => n11057, B2 => n10536, C1 => n11039, C2 =>
                           n10088, A => n8402, ZN => n8401);
   U15580 : OAI22_X1 port map( A1 => n580_port, A2 => n11584, B1 => n708_port, 
                           B2 => n11567, ZN => n8403);
   U15581 : AOI21_X1 port map( B1 => n8418, B2 => n8419, A => n10987, ZN => 
                           n8412);
   U15582 : AOI221_X1 port map( B1 => n11021, B2 => n10537, C1 => n11004, C2 =>
                           n10089, A => n8421, ZN => n8418);
   U15583 : AOI221_X1 port map( B1 => n11057, B2 => n10538, C1 => n11039, C2 =>
                           n10090, A => n8420, ZN => n8419);
   U15584 : OAI22_X1 port map( A1 => n579_port, A2 => n11584, B1 => n707_port, 
                           B2 => n11567, ZN => n8421);
   U15585 : AOI21_X1 port map( B1 => n8436, B2 => n8437, A => n10987, ZN => 
                           n8430);
   U15586 : AOI221_X1 port map( B1 => n11021, B2 => n10539, C1 => n11004, C2 =>
                           n10091, A => n8439, ZN => n8436);
   U15587 : AOI221_X1 port map( B1 => n11057, B2 => n10540, C1 => n11039, C2 =>
                           n10092, A => n8438, ZN => n8437);
   U15588 : OAI22_X1 port map( A1 => n578_port, A2 => n11584, B1 => n706_port, 
                           B2 => n11567, ZN => n8439);
   U15589 : AOI21_X1 port map( B1 => n8454, B2 => n8455, A => n10987, ZN => 
                           n8448);
   U15590 : AOI221_X1 port map( B1 => n11021, B2 => n10541, C1 => n11004, C2 =>
                           n10093, A => n8459, ZN => n8454);
   U15591 : AOI221_X1 port map( B1 => n11057, B2 => n10542, C1 => n11039, C2 =>
                           n10094, A => n8456, ZN => n8455);
   U15592 : OAI22_X1 port map( A1 => n577_port, A2 => n11584, B1 => n705_port, 
                           B2 => n11567, ZN => n8459);
   U15593 : AOI21_X1 port map( B1 => n8483, B2 => n8484, A => n10767, ZN => 
                           n8472);
   U15594 : AOI221_X1 port map( B1 => n10787, B2 => n10415, C1 => n10770, C2 =>
                           n9967, A => n8487, ZN => n8483);
   U15595 : AOI221_X1 port map( B1 => n10822, B2 => n10416, C1 => n10804, C2 =>
                           n9968, A => n8486, ZN => n8484);
   U15596 : OAI22_X1 port map( A1 => n640_port, A2 => n11662, B1 => n768_port, 
                           B2 => n11645, ZN => n8487);
   U15597 : AOI21_X1 port map( B1 => n8518, B2 => n8519, A => n10767, ZN => 
                           n8512);
   U15598 : AOI221_X1 port map( B1 => n10787, B2 => n10417, C1 => n10770, C2 =>
                           n9969, A => n8521, ZN => n8518);
   U15599 : AOI221_X1 port map( B1 => n10822, B2 => n10418, C1 => n10804, C2 =>
                           n9970, A => n8520, ZN => n8519);
   U15600 : OAI22_X1 port map( A1 => n639_port, A2 => n11662, B1 => n767_port, 
                           B2 => n11645, ZN => n8521);
   U15601 : AOI21_X1 port map( B1 => n8536, B2 => n8537, A => n10767, ZN => 
                           n8530);
   U15602 : AOI221_X1 port map( B1 => n10787, B2 => n10419, C1 => n10770, C2 =>
                           n9971, A => n8539, ZN => n8536);
   U15603 : AOI221_X1 port map( B1 => n10822, B2 => n10420, C1 => n10804, C2 =>
                           n9972, A => n8538, ZN => n8537);
   U15604 : OAI22_X1 port map( A1 => n638_port, A2 => n11662, B1 => n766_port, 
                           B2 => n11645, ZN => n8539);
   U15605 : AOI21_X1 port map( B1 => n8554, B2 => n8555, A => n10767, ZN => 
                           n8548);
   U15606 : AOI221_X1 port map( B1 => n10787, B2 => n10421, C1 => n10770, C2 =>
                           n9973, A => n8557, ZN => n8554);
   U15607 : AOI221_X1 port map( B1 => n10822, B2 => n10422, C1 => n10804, C2 =>
                           n9974, A => n8556, ZN => n8555);
   U15608 : OAI22_X1 port map( A1 => n637_port, A2 => n11662, B1 => n765_port, 
                           B2 => n11645, ZN => n8557);
   U15609 : AOI21_X1 port map( B1 => n8572, B2 => n8573, A => n10766, ZN => 
                           n8566);
   U15610 : AOI221_X1 port map( B1 => n10787, B2 => n10423, C1 => n10770, C2 =>
                           n9975, A => n8575, ZN => n8572);
   U15611 : AOI221_X1 port map( B1 => n10822, B2 => n10424, C1 => n10804, C2 =>
                           n9976, A => n8574, ZN => n8573);
   U15612 : OAI22_X1 port map( A1 => n636_port, A2 => n11661, B1 => n764_port, 
                           B2 => n11644, ZN => n8575);
   U15613 : AOI21_X1 port map( B1 => n8590, B2 => n8591, A => n10766, ZN => 
                           n8584);
   U15614 : AOI221_X1 port map( B1 => n10787, B2 => n10425, C1 => n10770, C2 =>
                           n9977, A => n8593, ZN => n8590);
   U15615 : AOI221_X1 port map( B1 => n10822, B2 => n10426, C1 => n10804, C2 =>
                           n9978, A => n8592, ZN => n8591);
   U15616 : OAI22_X1 port map( A1 => n635_port, A2 => n11661, B1 => n763_port, 
                           B2 => n11644, ZN => n8593);
   U15617 : AOI21_X1 port map( B1 => n8608, B2 => n8609, A => n10766, ZN => 
                           n8602);
   U15618 : AOI221_X1 port map( B1 => n10788, B2 => n10427, C1 => n10771, C2 =>
                           n9979, A => n8611, ZN => n8608);
   U15619 : AOI221_X1 port map( B1 => n10823, B2 => n10428, C1 => n10805, C2 =>
                           n9980, A => n8610, ZN => n8609);
   U15620 : OAI22_X1 port map( A1 => n634_port, A2 => n11661, B1 => n762_port, 
                           B2 => n11644, ZN => n8611);
   U15621 : AOI21_X1 port map( B1 => n8626, B2 => n8627, A => n10766, ZN => 
                           n8620);
   U15622 : AOI221_X1 port map( B1 => n10788, B2 => n10429, C1 => n10771, C2 =>
                           n9981, A => n8629, ZN => n8626);
   U15623 : AOI221_X1 port map( B1 => n10823, B2 => n10430, C1 => n10805, C2 =>
                           n9982, A => n8628, ZN => n8627);
   U15624 : OAI22_X1 port map( A1 => n633_port, A2 => n11661, B1 => n761_port, 
                           B2 => n11644, ZN => n8629);
   U15625 : AOI21_X1 port map( B1 => n8644, B2 => n8645, A => n10766, ZN => 
                           n8638);
   U15626 : AOI221_X1 port map( B1 => n10788, B2 => n10431, C1 => n10771, C2 =>
                           n9983, A => n8647, ZN => n8644);
   U15627 : AOI221_X1 port map( B1 => n10823, B2 => n10432, C1 => n10805, C2 =>
                           n9984, A => n8646, ZN => n8645);
   U15628 : OAI22_X1 port map( A1 => n632_port, A2 => n11661, B1 => n760_port, 
                           B2 => n11644, ZN => n8647);
   U15629 : AOI21_X1 port map( B1 => n8662, B2 => n8663, A => n10766, ZN => 
                           n8656);
   U15630 : AOI221_X1 port map( B1 => n10788, B2 => n10433, C1 => n10771, C2 =>
                           n9985, A => n8665, ZN => n8662);
   U15631 : AOI221_X1 port map( B1 => n10823, B2 => n10434, C1 => n10805, C2 =>
                           n9986, A => n8664, ZN => n8663);
   U15632 : OAI22_X1 port map( A1 => n631_port, A2 => n11661, B1 => n759_port, 
                           B2 => n11644, ZN => n8665);
   U15633 : AOI21_X1 port map( B1 => n8680, B2 => n8681, A => n10766, ZN => 
                           n8674);
   U15634 : AOI221_X1 port map( B1 => n10788, B2 => n10435, C1 => n10771, C2 =>
                           n9987, A => n8683, ZN => n8680);
   U15635 : AOI221_X1 port map( B1 => n10823, B2 => n10436, C1 => n10805, C2 =>
                           n9988, A => n8682, ZN => n8681);
   U15636 : OAI22_X1 port map( A1 => n630_port, A2 => n11660, B1 => n758_port, 
                           B2 => n11643, ZN => n8683);
   U15637 : AOI21_X1 port map( B1 => n8698, B2 => n8699, A => n10766, ZN => 
                           n8692);
   U15638 : AOI221_X1 port map( B1 => n10788, B2 => n10437, C1 => n10771, C2 =>
                           n9989, A => n8701, ZN => n8698);
   U15639 : AOI221_X1 port map( B1 => n10823, B2 => n10438, C1 => n10805, C2 =>
                           n9990, A => n8700, ZN => n8699);
   U15640 : OAI22_X1 port map( A1 => n629_port, A2 => n11660, B1 => n757_port, 
                           B2 => n11643, ZN => n8701);
   U15641 : AOI21_X1 port map( B1 => n8716, B2 => n8717, A => n10766, ZN => 
                           n8710);
   U15642 : AOI221_X1 port map( B1 => n10788, B2 => n10439, C1 => n10771, C2 =>
                           n9991, A => n8719, ZN => n8716);
   U15643 : AOI221_X1 port map( B1 => n10824, B2 => n10440, C1 => n10806, C2 =>
                           n9992, A => n8718, ZN => n8717);
   U15644 : OAI22_X1 port map( A1 => n628_port, A2 => n11660, B1 => n756_port, 
                           B2 => n11643, ZN => n8719);
   U15645 : AOI21_X1 port map( B1 => n8734, B2 => n8735, A => n10766, ZN => 
                           n8728);
   U15646 : AOI221_X1 port map( B1 => n10789, B2 => n10441, C1 => n10772, C2 =>
                           n9993, A => n8737, ZN => n8734);
   U15647 : AOI221_X1 port map( B1 => n10824, B2 => n10442, C1 => n10806, C2 =>
                           n9994, A => n8736, ZN => n8735);
   U15648 : OAI22_X1 port map( A1 => n627_port, A2 => n11660, B1 => n755_port, 
                           B2 => n11643, ZN => n8737);
   U15649 : AOI21_X1 port map( B1 => n8752, B2 => n8753, A => n10766, ZN => 
                           n8746);
   U15650 : AOI221_X1 port map( B1 => n10789, B2 => n10443, C1 => n10772, C2 =>
                           n9995, A => n8755, ZN => n8752);
   U15651 : AOI221_X1 port map( B1 => n10824, B2 => n10444, C1 => n10806, C2 =>
                           n9996, A => n8754, ZN => n8753);
   U15652 : OAI22_X1 port map( A1 => n626_port, A2 => n11660, B1 => n754_port, 
                           B2 => n11643, ZN => n8755);
   U15653 : AOI21_X1 port map( B1 => n8770, B2 => n8771, A => n10766, ZN => 
                           n8764);
   U15654 : AOI221_X1 port map( B1 => n10789, B2 => n10445, C1 => n10772, C2 =>
                           n9997, A => n8773, ZN => n8770);
   U15655 : AOI221_X1 port map( B1 => n10824, B2 => n10446, C1 => n10806, C2 =>
                           n9998, A => n8772, ZN => n8771);
   U15656 : OAI22_X1 port map( A1 => n625_port, A2 => n11660, B1 => n753_port, 
                           B2 => n11643, ZN => n8773);
   U15657 : AOI21_X1 port map( B1 => n8788, B2 => n8789, A => n10765, ZN => 
                           n8782);
   U15658 : AOI221_X1 port map( B1 => n10789, B2 => n10447, C1 => n10772, C2 =>
                           n9999, A => n8791, ZN => n8788);
   U15659 : AOI221_X1 port map( B1 => n10824, B2 => n10448, C1 => n10806, C2 =>
                           n10000, A => n8790, ZN => n8789);
   U15660 : OAI22_X1 port map( A1 => n624_port, A2 => n11659, B1 => n752_port, 
                           B2 => n11642, ZN => n8791);
   U15661 : AOI21_X1 port map( B1 => n8806, B2 => n8807, A => n10765, ZN => 
                           n8800);
   U15662 : AOI221_X1 port map( B1 => n10789, B2 => n10449, C1 => n10772, C2 =>
                           n10001, A => n8809, ZN => n8806);
   U15663 : AOI221_X1 port map( B1 => n10824, B2 => n10450, C1 => n10806, C2 =>
                           n10002, A => n8808, ZN => n8807);
   U15664 : OAI22_X1 port map( A1 => n623_port, A2 => n11659, B1 => n751_port, 
                           B2 => n11642, ZN => n8809);
   U15665 : AOI21_X1 port map( B1 => n8824, B2 => n8825, A => n10765, ZN => 
                           n8818);
   U15666 : AOI221_X1 port map( B1 => n10789, B2 => n10451, C1 => n10772, C2 =>
                           n10003, A => n8827, ZN => n8824);
   U15667 : AOI221_X1 port map( B1 => n10825, B2 => n10452, C1 => n10807, C2 =>
                           n10004, A => n8826, ZN => n8825);
   U15668 : OAI22_X1 port map( A1 => n622_port, A2 => n11659, B1 => n750_port, 
                           B2 => n11642, ZN => n8827);
   U15669 : AOI21_X1 port map( B1 => n8842, B2 => n8843, A => n10765, ZN => 
                           n8836);
   U15670 : AOI221_X1 port map( B1 => n10790, B2 => n10453, C1 => n10773, C2 =>
                           n10005, A => n8845, ZN => n8842);
   U15671 : AOI221_X1 port map( B1 => n10825, B2 => n10454, C1 => n10807, C2 =>
                           n10006, A => n8844, ZN => n8843);
   U15672 : OAI22_X1 port map( A1 => n621_port, A2 => n11659, B1 => n749_port, 
                           B2 => n11642, ZN => n8845);
   U15673 : AOI21_X1 port map( B1 => n8860, B2 => n8861, A => n10765, ZN => 
                           n8854);
   U15674 : AOI221_X1 port map( B1 => n10790, B2 => n10455, C1 => n10773, C2 =>
                           n10007, A => n8863, ZN => n8860);
   U15675 : AOI221_X1 port map( B1 => n10825, B2 => n10456, C1 => n10807, C2 =>
                           n10008, A => n8862, ZN => n8861);
   U15676 : OAI22_X1 port map( A1 => n620_port, A2 => n11659, B1 => n748_port, 
                           B2 => n11642, ZN => n8863);
   U15677 : AOI21_X1 port map( B1 => n8878, B2 => n8879, A => n10765, ZN => 
                           n8872);
   U15678 : AOI221_X1 port map( B1 => n10790, B2 => n10457, C1 => n10773, C2 =>
                           n10009, A => n8881, ZN => n8878);
   U15679 : AOI221_X1 port map( B1 => n10825, B2 => n10458, C1 => n10807, C2 =>
                           n10010, A => n8880, ZN => n8879);
   U15680 : OAI22_X1 port map( A1 => n619_port, A2 => n11659, B1 => n747_port, 
                           B2 => n11642, ZN => n8881);
   U15681 : AOI21_X1 port map( B1 => n8896, B2 => n8897, A => n10765, ZN => 
                           n8890);
   U15682 : AOI221_X1 port map( B1 => n10790, B2 => n10459, C1 => n10773, C2 =>
                           n10011, A => n8899, ZN => n8896);
   U15683 : AOI221_X1 port map( B1 => n10825, B2 => n10460, C1 => n10807, C2 =>
                           n10012, A => n8898, ZN => n8897);
   U15684 : OAI22_X1 port map( A1 => n618_port, A2 => n11658, B1 => n746_port, 
                           B2 => n11641, ZN => n8899);
   U15685 : AOI21_X1 port map( B1 => n8914, B2 => n8915, A => n10765, ZN => 
                           n8908);
   U15686 : AOI221_X1 port map( B1 => n10790, B2 => n10461, C1 => n10773, C2 =>
                           n10013, A => n8917, ZN => n8914);
   U15687 : AOI221_X1 port map( B1 => n10825, B2 => n10462, C1 => n10807, C2 =>
                           n10014, A => n8916, ZN => n8915);
   U15688 : OAI22_X1 port map( A1 => n617_port, A2 => n11658, B1 => n745_port, 
                           B2 => n11641, ZN => n8917);
   U15689 : AOI21_X1 port map( B1 => n8932, B2 => n8933, A => n10765, ZN => 
                           n8926);
   U15690 : AOI221_X1 port map( B1 => n10790, B2 => n10463, C1 => n10773, C2 =>
                           n10015, A => n8935, ZN => n8932);
   U15691 : AOI221_X1 port map( B1 => n10826, B2 => n10464, C1 => n10808, C2 =>
                           n10016, A => n8934, ZN => n8933);
   U15692 : OAI22_X1 port map( A1 => n616_port, A2 => n11658, B1 => n744_port, 
                           B2 => n11641, ZN => n8935);
   U15693 : AOI21_X1 port map( B1 => n8950, B2 => n8951, A => n10765, ZN => 
                           n8944);
   U15694 : AOI221_X1 port map( B1 => n10790, B2 => n10465, C1 => n10773, C2 =>
                           n10017, A => n8953, ZN => n8950);
   U15695 : AOI221_X1 port map( B1 => n10826, B2 => n10466, C1 => n10808, C2 =>
                           n10018, A => n8952, ZN => n8951);
   U15696 : OAI22_X1 port map( A1 => n615_port, A2 => n11658, B1 => n743_port, 
                           B2 => n11641, ZN => n8953);
   U15697 : AOI21_X1 port map( B1 => n8968, B2 => n8969, A => n10765, ZN => 
                           n8962);
   U15698 : AOI221_X1 port map( B1 => n10791, B2 => n10467, C1 => n10774, C2 =>
                           n10019, A => n8971, ZN => n8968);
   U15699 : AOI221_X1 port map( B1 => n10826, B2 => n10468, C1 => n10808, C2 =>
                           n10020, A => n8970, ZN => n8969);
   U15700 : OAI22_X1 port map( A1 => n614_port, A2 => n11658, B1 => n742_port, 
                           B2 => n11641, ZN => n8971);
   U15701 : AOI21_X1 port map( B1 => n8986, B2 => n8987, A => n10765, ZN => 
                           n8980);
   U15702 : AOI221_X1 port map( B1 => n10791, B2 => n10469, C1 => n10774, C2 =>
                           n10021, A => n8989, ZN => n8986);
   U15703 : AOI221_X1 port map( B1 => n10826, B2 => n10470, C1 => n10808, C2 =>
                           n10022, A => n8988, ZN => n8987);
   U15704 : OAI22_X1 port map( A1 => n613_port, A2 => n11658, B1 => n741_port, 
                           B2 => n11641, ZN => n8989);
   U15705 : AOI21_X1 port map( B1 => n9004, B2 => n9005, A => n10764, ZN => 
                           n8998);
   U15706 : AOI221_X1 port map( B1 => n10791, B2 => n10471, C1 => n10774, C2 =>
                           n10023, A => n9007, ZN => n9004);
   U15707 : AOI221_X1 port map( B1 => n10826, B2 => n10472, C1 => n10808, C2 =>
                           n10024, A => n9006, ZN => n9005);
   U15708 : OAI22_X1 port map( A1 => n612_port, A2 => n11657, B1 => n740_port, 
                           B2 => n11640, ZN => n9007);
   U15709 : AOI21_X1 port map( B1 => n9022, B2 => n9023, A => n10764, ZN => 
                           n9016);
   U15710 : AOI221_X1 port map( B1 => n10791, B2 => n10473, C1 => n10774, C2 =>
                           n10025, A => n9025, ZN => n9022);
   U15711 : AOI221_X1 port map( B1 => n10826, B2 => n10474, C1 => n10808, C2 =>
                           n10026, A => n9024, ZN => n9023);
   U15712 : OAI22_X1 port map( A1 => n611_port, A2 => n11657, B1 => n739_port, 
                           B2 => n11640, ZN => n9025);
   U15713 : AOI21_X1 port map( B1 => n9040, B2 => n9041, A => n10764, ZN => 
                           n9034);
   U15714 : AOI221_X1 port map( B1 => n10791, B2 => n10475, C1 => n10774, C2 =>
                           n10027, A => n9043, ZN => n9040);
   U15715 : AOI221_X1 port map( B1 => n10827, B2 => n10476, C1 => n10809, C2 =>
                           n10028, A => n9042, ZN => n9041);
   U15716 : OAI22_X1 port map( A1 => n610_port, A2 => n11657, B1 => n738_port, 
                           B2 => n11640, ZN => n9043);
   U15717 : AOI21_X1 port map( B1 => n9058, B2 => n9059, A => n10764, ZN => 
                           n9052);
   U15718 : AOI221_X1 port map( B1 => n10791, B2 => n10477, C1 => n10774, C2 =>
                           n10029, A => n9061, ZN => n9058);
   U15719 : AOI221_X1 port map( B1 => n10827, B2 => n10478, C1 => n10809, C2 =>
                           n10030, A => n9060, ZN => n9059);
   U15720 : OAI22_X1 port map( A1 => n609_port, A2 => n11657, B1 => n737_port, 
                           B2 => n11640, ZN => n9061);
   U15721 : AOI21_X1 port map( B1 => n9076, B2 => n9077, A => n10764, ZN => 
                           n9070);
   U15722 : AOI221_X1 port map( B1 => n10792, B2 => n10479, C1 => n10775, C2 =>
                           n10031, A => n9079, ZN => n9076);
   U15723 : AOI221_X1 port map( B1 => n10827, B2 => n10480, C1 => n10809, C2 =>
                           n10032, A => n9078, ZN => n9077);
   U15724 : OAI22_X1 port map( A1 => n608_port, A2 => n11657, B1 => n736_port, 
                           B2 => n11640, ZN => n9079);
   U15725 : AOI21_X1 port map( B1 => n9094, B2 => n9095, A => n10764, ZN => 
                           n9088);
   U15726 : AOI221_X1 port map( B1 => n10792, B2 => n10481, C1 => n10775, C2 =>
                           n10033, A => n9097, ZN => n9094);
   U15727 : AOI221_X1 port map( B1 => n10827, B2 => n10482, C1 => n10809, C2 =>
                           n10034, A => n9096, ZN => n9095);
   U15728 : OAI22_X1 port map( A1 => n607_port, A2 => n11657, B1 => n735_port, 
                           B2 => n11640, ZN => n9097);
   U15729 : AOI21_X1 port map( B1 => n9112, B2 => n9113, A => n10764, ZN => 
                           n9106);
   U15730 : AOI221_X1 port map( B1 => n10792, B2 => n10483, C1 => n10775, C2 =>
                           n10035, A => n9115, ZN => n9112);
   U15731 : AOI221_X1 port map( B1 => n10827, B2 => n10484, C1 => n10809, C2 =>
                           n10036, A => n9114, ZN => n9113);
   U15732 : OAI22_X1 port map( A1 => n606_port, A2 => n11656, B1 => n734_port, 
                           B2 => n11639, ZN => n9115);
   U15733 : AOI21_X1 port map( B1 => n9130, B2 => n9131, A => n10764, ZN => 
                           n9124);
   U15734 : AOI221_X1 port map( B1 => n10792, B2 => n10485, C1 => n10775, C2 =>
                           n10037, A => n9133, ZN => n9130);
   U15735 : AOI221_X1 port map( B1 => n10827, B2 => n10486, C1 => n10809, C2 =>
                           n10038, A => n9132, ZN => n9131);
   U15736 : OAI22_X1 port map( A1 => n605_port, A2 => n11656, B1 => n733_port, 
                           B2 => n11639, ZN => n9133);
   U15737 : AOI21_X1 port map( B1 => n9148, B2 => n9149, A => n10764, ZN => 
                           n9142);
   U15738 : AOI221_X1 port map( B1 => n10792, B2 => n10487, C1 => n10775, C2 =>
                           n10039, A => n9151, ZN => n9148);
   U15739 : AOI221_X1 port map( B1 => n10828, B2 => n10488, C1 => n10810, C2 =>
                           n10040, A => n9150, ZN => n9149);
   U15740 : OAI22_X1 port map( A1 => n604_port, A2 => n11656, B1 => n732_port, 
                           B2 => n11639, ZN => n9151);
   U15741 : AOI21_X1 port map( B1 => n9166, B2 => n9167, A => n10764, ZN => 
                           n9160);
   U15742 : AOI221_X1 port map( B1 => n10792, B2 => n10489, C1 => n10775, C2 =>
                           n10041, A => n9169, ZN => n9166);
   U15743 : AOI221_X1 port map( B1 => n10828, B2 => n10490, C1 => n10810, C2 =>
                           n10042, A => n9168, ZN => n9167);
   U15744 : OAI22_X1 port map( A1 => n603_port, A2 => n11656, B1 => n731_port, 
                           B2 => n11639, ZN => n9169);
   U15745 : AOI21_X1 port map( B1 => n9184, B2 => n9185, A => n10764, ZN => 
                           n9178);
   U15746 : AOI221_X1 port map( B1 => n10793, B2 => n10491, C1 => n10776, C2 =>
                           n10043, A => n9187, ZN => n9184);
   U15747 : AOI221_X1 port map( B1 => n10828, B2 => n10492, C1 => n10810, C2 =>
                           n10044, A => n9186, ZN => n9185);
   U15748 : OAI22_X1 port map( A1 => n602_port, A2 => n11656, B1 => n730_port, 
                           B2 => n11639, ZN => n9187);
   U15749 : AOI21_X1 port map( B1 => n9202, B2 => n9203, A => n10764, ZN => 
                           n9196);
   U15750 : AOI221_X1 port map( B1 => n10793, B2 => n10493, C1 => n10776, C2 =>
                           n10045, A => n9205, ZN => n9202);
   U15751 : AOI221_X1 port map( B1 => n10828, B2 => n10494, C1 => n10810, C2 =>
                           n10046, A => n9204, ZN => n9203);
   U15752 : OAI22_X1 port map( A1 => n601_port, A2 => n11656, B1 => n729_port, 
                           B2 => n11639, ZN => n9205);
   U15753 : AOI21_X1 port map( B1 => n9220, B2 => n9221, A => n10763, ZN => 
                           n9214);
   U15754 : AOI221_X1 port map( B1 => n10793, B2 => n10495, C1 => n10776, C2 =>
                           n10047, A => n9223, ZN => n9220);
   U15755 : AOI221_X1 port map( B1 => n10828, B2 => n10496, C1 => n10810, C2 =>
                           n10048, A => n9222, ZN => n9221);
   U15756 : OAI22_X1 port map( A1 => n600_port, A2 => n11655, B1 => n728_port, 
                           B2 => n11638, ZN => n9223);
   U15757 : AOI21_X1 port map( B1 => n9238, B2 => n9239, A => n10763, ZN => 
                           n9232);
   U15758 : AOI221_X1 port map( B1 => n10793, B2 => n10497, C1 => n10776, C2 =>
                           n10049, A => n9241, ZN => n9238);
   U15759 : AOI221_X1 port map( B1 => n10828, B2 => n10498, C1 => n10810, C2 =>
                           n10050, A => n9240, ZN => n9239);
   U15760 : OAI22_X1 port map( A1 => n599_port, A2 => n11655, B1 => n727_port, 
                           B2 => n11638, ZN => n9241);
   U15761 : AOI21_X1 port map( B1 => n9256, B2 => n9257, A => n10763, ZN => 
                           n9250);
   U15762 : AOI221_X1 port map( B1 => n10793, B2 => n10499, C1 => n10776, C2 =>
                           n10051, A => n9259, ZN => n9256);
   U15763 : AOI221_X1 port map( B1 => n10829, B2 => n10500, C1 => n10811, C2 =>
                           n10052, A => n9258, ZN => n9257);
   U15764 : OAI22_X1 port map( A1 => n598_port, A2 => n11655, B1 => n726_port, 
                           B2 => n11638, ZN => n9259);
   U15765 : AOI21_X1 port map( B1 => n9274, B2 => n9275, A => n10763, ZN => 
                           n9268);
   U15766 : AOI221_X1 port map( B1 => n10793, B2 => n10501, C1 => n10776, C2 =>
                           n10053, A => n9277, ZN => n9274);
   U15767 : AOI221_X1 port map( B1 => n10829, B2 => n10502, C1 => n10811, C2 =>
                           n10054, A => n9276, ZN => n9275);
   U15768 : OAI22_X1 port map( A1 => n597_port, A2 => n11655, B1 => n725_port, 
                           B2 => n11638, ZN => n9277);
   U15769 : AOI21_X1 port map( B1 => n9292, B2 => n9293, A => n10763, ZN => 
                           n9286);
   U15770 : AOI221_X1 port map( B1 => n10793, B2 => n10503, C1 => n10776, C2 =>
                           n10055, A => n9295, ZN => n9292);
   U15771 : AOI221_X1 port map( B1 => n10829, B2 => n10504, C1 => n10811, C2 =>
                           n10056, A => n9294, ZN => n9293);
   U15772 : OAI22_X1 port map( A1 => n596_port, A2 => n11655, B1 => n724_port, 
                           B2 => n11638, ZN => n9295);
   U15773 : AOI21_X1 port map( B1 => n9310, B2 => n9311, A => n10763, ZN => 
                           n9304);
   U15774 : AOI221_X1 port map( B1 => n10794, B2 => n10505, C1 => n10777, C2 =>
                           n10057, A => n9313, ZN => n9310);
   U15775 : AOI221_X1 port map( B1 => n10829, B2 => n10506, C1 => n10811, C2 =>
                           n10058, A => n9312, ZN => n9311);
   U15776 : OAI22_X1 port map( A1 => n595_port, A2 => n11655, B1 => n723_port, 
                           B2 => n11638, ZN => n9313);
   U15777 : AOI21_X1 port map( B1 => n9328, B2 => n9329, A => n10763, ZN => 
                           n9322);
   U15778 : AOI221_X1 port map( B1 => n10794, B2 => n10507, C1 => n10777, C2 =>
                           n10059, A => n9331, ZN => n9328);
   U15779 : AOI221_X1 port map( B1 => n10829, B2 => n10508, C1 => n10811, C2 =>
                           n10060, A => n9330, ZN => n9329);
   U15780 : OAI22_X1 port map( A1 => n594_port, A2 => n11654, B1 => n722_port, 
                           B2 => n11637, ZN => n9331);
   U15781 : AOI21_X1 port map( B1 => n9346, B2 => n9347, A => n10763, ZN => 
                           n9340);
   U15782 : AOI221_X1 port map( B1 => n10794, B2 => n10509, C1 => n10777, C2 =>
                           n10061, A => n9349, ZN => n9346);
   U15783 : AOI221_X1 port map( B1 => n10829, B2 => n10510, C1 => n10811, C2 =>
                           n10062, A => n9348, ZN => n9347);
   U15784 : OAI22_X1 port map( A1 => n593_port, A2 => n11654, B1 => n721_port, 
                           B2 => n11637, ZN => n9349);
   U15785 : AOI21_X1 port map( B1 => n9364, B2 => n9365, A => n10763, ZN => 
                           n9358);
   U15786 : AOI221_X1 port map( B1 => n10794, B2 => n10511, C1 => n10777, C2 =>
                           n10063, A => n9367, ZN => n9364);
   U15787 : AOI221_X1 port map( B1 => n10830, B2 => n10512, C1 => n10812, C2 =>
                           n10064, A => n9366, ZN => n9365);
   U15788 : OAI22_X1 port map( A1 => n592_port, A2 => n11654, B1 => n720_port, 
                           B2 => n11637, ZN => n9367);
   U15789 : AOI21_X1 port map( B1 => n9382, B2 => n9383, A => n10763, ZN => 
                           n9376);
   U15790 : AOI221_X1 port map( B1 => n10794, B2 => n10513, C1 => n10777, C2 =>
                           n10065, A => n9385, ZN => n9382);
   U15791 : AOI221_X1 port map( B1 => n10830, B2 => n10514, C1 => n10812, C2 =>
                           n10066, A => n9384, ZN => n9383);
   U15792 : OAI22_X1 port map( A1 => n591_port, A2 => n11654, B1 => n719_port, 
                           B2 => n11637, ZN => n9385);
   U15793 : AOI21_X1 port map( B1 => n9400, B2 => n9401, A => n10763, ZN => 
                           n9394);
   U15794 : AOI221_X1 port map( B1 => n10794, B2 => n10515, C1 => n10777, C2 =>
                           n10067, A => n9403, ZN => n9400);
   U15795 : AOI221_X1 port map( B1 => n10830, B2 => n10516, C1 => n10812, C2 =>
                           n10068, A => n9402, ZN => n9401);
   U15796 : OAI22_X1 port map( A1 => n590_port, A2 => n11654, B1 => n718_port, 
                           B2 => n11637, ZN => n9403);
   U15797 : AOI21_X1 port map( B1 => n9418, B2 => n9419, A => n10763, ZN => 
                           n9412);
   U15798 : AOI221_X1 port map( B1 => n10795, B2 => n10517, C1 => n10778, C2 =>
                           n10069, A => n9421, ZN => n9418);
   U15799 : AOI221_X1 port map( B1 => n10830, B2 => n10518, C1 => n10812, C2 =>
                           n10070, A => n9420, ZN => n9419);
   U15800 : OAI22_X1 port map( A1 => n589_port, A2 => n11654, B1 => n717_port, 
                           B2 => n11637, ZN => n9421);
   U15801 : AOI21_X1 port map( B1 => n9436, B2 => n9437, A => n10762, ZN => 
                           n9430);
   U15802 : AOI221_X1 port map( B1 => n10795, B2 => n10519, C1 => n10778, C2 =>
                           n10071, A => n9439, ZN => n9436);
   U15803 : AOI221_X1 port map( B1 => n10830, B2 => n10520, C1 => n10812, C2 =>
                           n10072, A => n9438, ZN => n9437);
   U15804 : OAI22_X1 port map( A1 => n588_port, A2 => n11653, B1 => n716_port, 
                           B2 => n11636, ZN => n9439);
   U15805 : AOI21_X1 port map( B1 => n9454, B2 => n9455, A => n10762, ZN => 
                           n9448);
   U15806 : AOI221_X1 port map( B1 => n10795, B2 => n10521, C1 => n10778, C2 =>
                           n10073, A => n9457, ZN => n9454);
   U15807 : AOI221_X1 port map( B1 => n10830, B2 => n10522, C1 => n10812, C2 =>
                           n10074, A => n9456, ZN => n9455);
   U15808 : OAI22_X1 port map( A1 => n587_port, A2 => n11653, B1 => n715_port, 
                           B2 => n11636, ZN => n9457);
   U15809 : AOI21_X1 port map( B1 => n9472, B2 => n9473, A => n10762, ZN => 
                           n9466);
   U15810 : AOI221_X1 port map( B1 => n10795, B2 => n10523, C1 => n10778, C2 =>
                           n10075, A => n9475, ZN => n9472);
   U15811 : AOI221_X1 port map( B1 => n10831, B2 => n10524, C1 => n10813, C2 =>
                           n10076, A => n9474, ZN => n9473);
   U15812 : OAI22_X1 port map( A1 => n586_port, A2 => n11653, B1 => n714_port, 
                           B2 => n11636, ZN => n9475);
   U15813 : AOI21_X1 port map( B1 => n9490, B2 => n9491, A => n10762, ZN => 
                           n9484);
   U15814 : AOI221_X1 port map( B1 => n10795, B2 => n10525, C1 => n10778, C2 =>
                           n10077, A => n9493, ZN => n9490);
   U15815 : AOI221_X1 port map( B1 => n10831, B2 => n10526, C1 => n10813, C2 =>
                           n10078, A => n9492, ZN => n9491);
   U15816 : OAI22_X1 port map( A1 => n585_port, A2 => n11653, B1 => n713_port, 
                           B2 => n11636, ZN => n9493);
   U15817 : AOI21_X1 port map( B1 => n9508, B2 => n9509, A => n10762, ZN => 
                           n9502);
   U15818 : AOI221_X1 port map( B1 => n10795, B2 => n10527, C1 => n10778, C2 =>
                           n10079, A => n9511, ZN => n9508);
   U15819 : AOI221_X1 port map( B1 => n10831, B2 => n10528, C1 => n10813, C2 =>
                           n10080, A => n9510, ZN => n9509);
   U15820 : OAI22_X1 port map( A1 => n584_port, A2 => n11653, B1 => n712_port, 
                           B2 => n11636, ZN => n9511);
   U15821 : AOI21_X1 port map( B1 => n9526, B2 => n9527, A => n10762, ZN => 
                           n9520);
   U15822 : AOI221_X1 port map( B1 => n10795, B2 => n10529, C1 => n10778, C2 =>
                           n10081, A => n9529, ZN => n9526);
   U15823 : AOI221_X1 port map( B1 => n10831, B2 => n10530, C1 => n10813, C2 =>
                           n10082, A => n9528, ZN => n9527);
   U15824 : OAI22_X1 port map( A1 => n583_port, A2 => n11653, B1 => n711_port, 
                           B2 => n11636, ZN => n9529);
   U15825 : AOI21_X1 port map( B1 => n9544, B2 => n9545, A => n10762, ZN => 
                           n9538);
   U15826 : AOI221_X1 port map( B1 => n10796, B2 => n10531, C1 => n10779, C2 =>
                           n10083, A => n9547, ZN => n9544);
   U15827 : AOI221_X1 port map( B1 => n10831, B2 => n10532, C1 => n10813, C2 =>
                           n10084, A => n9546, ZN => n9545);
   U15828 : OAI22_X1 port map( A1 => n582_port, A2 => n11652, B1 => n710_port, 
                           B2 => n11635, ZN => n9547);
   U15829 : AOI21_X1 port map( B1 => n9562, B2 => n9563, A => n10762, ZN => 
                           n9556);
   U15830 : AOI221_X1 port map( B1 => n10796, B2 => n10533, C1 => n10779, C2 =>
                           n10085, A => n9565, ZN => n9562);
   U15831 : AOI221_X1 port map( B1 => n10831, B2 => n10534, C1 => n10813, C2 =>
                           n10086, A => n9564, ZN => n9563);
   U15832 : OAI22_X1 port map( A1 => n581_port, A2 => n11652, B1 => n709_port, 
                           B2 => n11635, ZN => n9565);
   U15833 : AOI21_X1 port map( B1 => n9580, B2 => n9581, A => n10762, ZN => 
                           n9574);
   U15834 : AOI221_X1 port map( B1 => n10796, B2 => n10535, C1 => n10779, C2 =>
                           n10087, A => n9583, ZN => n9580);
   U15835 : AOI221_X1 port map( B1 => n10832, B2 => n10536, C1 => n10814, C2 =>
                           n10088, A => n9582, ZN => n9581);
   U15836 : OAI22_X1 port map( A1 => n580_port, A2 => n11652, B1 => n708_port, 
                           B2 => n11635, ZN => n9583);
   U15837 : AOI21_X1 port map( B1 => n9598, B2 => n9599, A => n10762, ZN => 
                           n9592);
   U15838 : AOI221_X1 port map( B1 => n10796, B2 => n10537, C1 => n10779, C2 =>
                           n10089, A => n9601, ZN => n9598);
   U15839 : AOI221_X1 port map( B1 => n10832, B2 => n10538, C1 => n10814, C2 =>
                           n10090, A => n9600, ZN => n9599);
   U15840 : OAI22_X1 port map( A1 => n579_port, A2 => n11652, B1 => n707_port, 
                           B2 => n11635, ZN => n9601);
   U15841 : AOI21_X1 port map( B1 => n9616, B2 => n9617, A => n10762, ZN => 
                           n9610);
   U15842 : AOI221_X1 port map( B1 => n10796, B2 => n10539, C1 => n10779, C2 =>
                           n10091, A => n9619, ZN => n9616);
   U15843 : AOI221_X1 port map( B1 => n10832, B2 => n10540, C1 => n10814, C2 =>
                           n10092, A => n9618, ZN => n9617);
   U15844 : OAI22_X1 port map( A1 => n578_port, A2 => n11652, B1 => n706_port, 
                           B2 => n11635, ZN => n9619);
   U15845 : AOI21_X1 port map( B1 => n9634, B2 => n9635, A => n10762, ZN => 
                           n9628);
   U15846 : AOI221_X1 port map( B1 => n10796, B2 => n10541, C1 => n10779, C2 =>
                           n10093, A => n9639, ZN => n9634);
   U15847 : AOI221_X1 port map( B1 => n10832, B2 => n10542, C1 => n10814, C2 =>
                           n10094, A => n9636, ZN => n9635);
   U15848 : OAI22_X1 port map( A1 => n577_port, A2 => n11652, B1 => n705_port, 
                           B2 => n11635, ZN => n9639);
   U15849 : INV_X1 port map( A => ADD_RD2(2), ZN => n6247);
   U15850 : INV_X1 port map( A => ADD_RD1(2), ZN => n6238);
   U15851 : INV_X1 port map( A => ADD_RD2(1), ZN => n6248);
   U15852 : INV_X1 port map( A => ADD_RD1(1), ZN => n6239);
   U15853 : INV_X1 port map( A => ADD_RD2(0), ZN => n6249);
   U15854 : INV_X1 port map( A => ADD_RD1(0), ZN => n6240);
   U15855 : INV_X1 port map( A => ADD_RD2(4), ZN => n6241);
   U15856 : INV_X1 port map( A => ADD_RD1(4), ZN => n6232);
   U15857 : OAI21_X1 port map( B1 => n2048_port, B2 => n11453, A => n11075, ZN 
                           => N2235);
   U15858 : OAI21_X1 port map( B1 => n2047_port, B2 => n11453, A => n11079, ZN 
                           => N2236);
   U15859 : OAI21_X1 port map( B1 => n2046_port, B2 => n11453, A => n11083, ZN 
                           => N2237);
   U15860 : OAI21_X1 port map( B1 => n2045_port, B2 => n11453, A => n11087, ZN 
                           => N2238);
   U15861 : OAI21_X1 port map( B1 => n2044_port, B2 => n11453, A => n11091, ZN 
                           => N2239);
   U15862 : OAI21_X1 port map( B1 => n2043_port, B2 => n11453, A => n11095, ZN 
                           => N2240);
   U15863 : OAI21_X1 port map( B1 => n2042_port, B2 => n11453, A => n11099, ZN 
                           => N2241);
   U15864 : OAI21_X1 port map( B1 => n2041_port, B2 => n11452, A => n11103, ZN 
                           => N2242);
   U15865 : OAI21_X1 port map( B1 => n2040_port, B2 => n11452, A => n11107, ZN 
                           => N2243);
   U15866 : OAI21_X1 port map( B1 => n2039_port, B2 => n11452, A => n11111, ZN 
                           => N2244);
   U15867 : OAI21_X1 port map( B1 => n2038_port, B2 => n11452, A => n11115, ZN 
                           => N2245);
   U15868 : OAI21_X1 port map( B1 => n2037_port, B2 => n11452, A => n11119, ZN 
                           => N2246);
   U15869 : OAI21_X1 port map( B1 => n2036_port, B2 => n11452, A => n11123, ZN 
                           => N2247);
   U15870 : OAI21_X1 port map( B1 => n2035_port, B2 => n11452, A => n11127, ZN 
                           => N2248);
   U15871 : OAI21_X1 port map( B1 => n2034_port, B2 => n11452, A => n11131, ZN 
                           => N2249);
   U15872 : OAI21_X1 port map( B1 => n2033_port, B2 => n11452, A => n11135, ZN 
                           => N2250);
   U15873 : OAI21_X1 port map( B1 => n2032_port, B2 => n11452, A => n11139, ZN 
                           => N2251);
   U15874 : OAI21_X1 port map( B1 => n2031_port, B2 => n11452, A => n11143, ZN 
                           => N2252);
   U15875 : OAI21_X1 port map( B1 => n2030_port, B2 => n11452, A => n11147, ZN 
                           => N2253);
   U15876 : OAI21_X1 port map( B1 => n2029_port, B2 => n11451, A => n11151, ZN 
                           => N2254);
   U15877 : OAI21_X1 port map( B1 => n2028_port, B2 => n11451, A => n11155, ZN 
                           => N2255);
   U15878 : OAI21_X1 port map( B1 => n2027_port, B2 => n11451, A => n11159, ZN 
                           => N2256);
   U15879 : OAI21_X1 port map( B1 => n2026_port, B2 => n11451, A => n11163, ZN 
                           => N2257);
   U15880 : OAI21_X1 port map( B1 => n2025_port, B2 => n11451, A => n11167, ZN 
                           => N2258);
   U15881 : OAI21_X1 port map( B1 => n2024_port, B2 => n11451, A => n11171, ZN 
                           => N2259);
   U15882 : OAI21_X1 port map( B1 => n2023_port, B2 => n11451, A => n11175, ZN 
                           => N2260);
   U15883 : OAI21_X1 port map( B1 => n2022_port, B2 => n11451, A => n11179, ZN 
                           => N2261);
   U15884 : OAI21_X1 port map( B1 => n2021_port, B2 => n11451, A => n11183, ZN 
                           => N2262);
   U15885 : OAI21_X1 port map( B1 => n2020_port, B2 => n11451, A => n11187, ZN 
                           => N2263);
   U15886 : OAI21_X1 port map( B1 => n2019_port, B2 => n11451, A => n11191, ZN 
                           => N2264);
   U15887 : OAI21_X1 port map( B1 => n2018_port, B2 => n11451, A => n11195, ZN 
                           => N2265);
   U15888 : OAI21_X1 port map( B1 => n2017_port, B2 => n11450, A => n11199, ZN 
                           => N2266);
   U15889 : OAI21_X1 port map( B1 => n2016_port, B2 => n11450, A => n11203, ZN 
                           => N2267);
   U15890 : OAI21_X1 port map( B1 => n2015_port, B2 => n11450, A => n11207, ZN 
                           => N2268);
   U15891 : OAI21_X1 port map( B1 => n2014_port, B2 => n11450, A => n11211, ZN 
                           => N2269);
   U15892 : OAI21_X1 port map( B1 => n2013_port, B2 => n11450, A => n11215, ZN 
                           => N2270);
   U15893 : OAI21_X1 port map( B1 => n2012_port, B2 => n11450, A => n11219, ZN 
                           => N2271);
   U15894 : OAI21_X1 port map( B1 => n2011_port, B2 => n11450, A => n11223, ZN 
                           => N2272);
   U15895 : OAI21_X1 port map( B1 => n2010_port, B2 => n11450, A => n11227, ZN 
                           => N2273);
   U15896 : OAI21_X1 port map( B1 => n2009_port, B2 => n11450, A => n11231, ZN 
                           => N2274);
   U15897 : OAI21_X1 port map( B1 => n2008_port, B2 => n11450, A => n11235, ZN 
                           => N2275);
   U15898 : OAI21_X1 port map( B1 => n2007_port, B2 => n11450, A => n11239, ZN 
                           => N2276);
   U15899 : OAI21_X1 port map( B1 => n2006_port, B2 => n11450, A => n11243, ZN 
                           => N2277);
   U15900 : OAI21_X1 port map( B1 => n2005_port, B2 => n11449, A => n11247, ZN 
                           => N2278);
   U15901 : OAI21_X1 port map( B1 => n2004_port, B2 => n11449, A => n11251, ZN 
                           => N2279);
   U15902 : OAI21_X1 port map( B1 => n2003_port, B2 => n11449, A => n11255, ZN 
                           => N2280);
   U15903 : OAI21_X1 port map( B1 => n2002_port, B2 => n11449, A => n11259, ZN 
                           => N2281);
   U15904 : OAI21_X1 port map( B1 => n2001_port, B2 => n11449, A => n11263, ZN 
                           => N2282);
   U15905 : OAI21_X1 port map( B1 => n2000_port, B2 => n11449, A => n11267, ZN 
                           => N2283);
   U15906 : OAI21_X1 port map( B1 => n1999_port, B2 => n11449, A => n11271, ZN 
                           => N2284);
   U15907 : OAI21_X1 port map( B1 => n1998_port, B2 => n11449, A => n11275, ZN 
                           => N2285);
   U15908 : OAI21_X1 port map( B1 => n1997_port, B2 => n11449, A => n11279, ZN 
                           => N2286);
   U15909 : OAI21_X1 port map( B1 => n1996_port, B2 => n11449, A => n11283, ZN 
                           => N2287);
   U15910 : OAI21_X1 port map( B1 => n1995_port, B2 => n11449, A => n11287, ZN 
                           => N2288);
   U15911 : OAI21_X1 port map( B1 => n1994_port, B2 => n11449, A => n11291, ZN 
                           => N2289);
   U15912 : OAI21_X1 port map( B1 => n1993_port, B2 => n11448, A => n11295, ZN 
                           => N2290);
   U15913 : OAI21_X1 port map( B1 => n1992_port, B2 => n11448, A => n11299, ZN 
                           => N2291);
   U15914 : OAI21_X1 port map( B1 => n1991_port, B2 => n11448, A => n11303, ZN 
                           => N2292);
   U15915 : OAI21_X1 port map( B1 => n1990_port, B2 => n11448, A => n11307, ZN 
                           => N2293);
   U15916 : OAI21_X1 port map( B1 => n1989_port, B2 => n11448, A => n11311, ZN 
                           => N2294);
   U15917 : OAI21_X1 port map( B1 => n1988_port, B2 => n11448, A => n11315, ZN 
                           => N2295);
   U15918 : OAI21_X1 port map( B1 => n1987_port, B2 => n11448, A => n11319, ZN 
                           => N2296);
   U15919 : OAI21_X1 port map( B1 => n1986_port, B2 => n11448, A => n11323, ZN 
                           => N2297);
   U15920 : OAI21_X1 port map( B1 => n1985_port, B2 => n11448, A => n11327, ZN 
                           => N2298);
   U15921 : OAI21_X1 port map( B1 => n1984_port, B2 => n11448, A => n11075, ZN 
                           => N2300);
   U15922 : OAI21_X1 port map( B1 => n1983_port, B2 => n11448, A => n11079, ZN 
                           => N2301);
   U15923 : OAI21_X1 port map( B1 => n1982_port, B2 => n11447, A => n11083, ZN 
                           => N2302);
   U15924 : OAI21_X1 port map( B1 => n1981_port, B2 => n11447, A => n11087, ZN 
                           => N2303);
   U15925 : OAI21_X1 port map( B1 => n1980_port, B2 => n11447, A => n11091, ZN 
                           => N2304);
   U15926 : OAI21_X1 port map( B1 => n1979_port, B2 => n11447, A => n11095, ZN 
                           => N2305);
   U15927 : OAI21_X1 port map( B1 => n1978_port, B2 => n11447, A => n11099, ZN 
                           => N2306);
   U15928 : OAI21_X1 port map( B1 => n1977_port, B2 => n11447, A => n11103, ZN 
                           => N2307);
   U15929 : OAI21_X1 port map( B1 => n1976_port, B2 => n11447, A => n11107, ZN 
                           => N2308);
   U15930 : OAI21_X1 port map( B1 => n1975_port, B2 => n11447, A => n11111, ZN 
                           => N2309);
   U15931 : OAI21_X1 port map( B1 => n1974_port, B2 => n11447, A => n11115, ZN 
                           => N2310);
   U15932 : OAI21_X1 port map( B1 => n1973_port, B2 => n11447, A => n11119, ZN 
                           => N2311);
   U15933 : OAI21_X1 port map( B1 => n1972_port, B2 => n11447, A => n11123, ZN 
                           => N2312);
   U15934 : OAI21_X1 port map( B1 => n1971_port, B2 => n11447, A => n11127, ZN 
                           => N2313);
   U15935 : OAI21_X1 port map( B1 => n1970_port, B2 => n11446, A => n11131, ZN 
                           => N2314);
   U15936 : OAI21_X1 port map( B1 => n1969_port, B2 => n11446, A => n11135, ZN 
                           => N2315);
   U15937 : OAI21_X1 port map( B1 => n1968_port, B2 => n11446, A => n11139, ZN 
                           => N2316);
   U15938 : OAI21_X1 port map( B1 => n1967_port, B2 => n11446, A => n11143, ZN 
                           => N2317);
   U15939 : OAI21_X1 port map( B1 => n1966_port, B2 => n11446, A => n11147, ZN 
                           => N2318);
   U15940 : OAI21_X1 port map( B1 => n1965_port, B2 => n11446, A => n11151, ZN 
                           => N2319);
   U15941 : OAI21_X1 port map( B1 => n1964_port, B2 => n11446, A => n11155, ZN 
                           => N2320);
   U15942 : OAI21_X1 port map( B1 => n1963_port, B2 => n11446, A => n11159, ZN 
                           => N2321);
   U15943 : OAI21_X1 port map( B1 => n1962_port, B2 => n11446, A => n11163, ZN 
                           => N2322);
   U15944 : OAI21_X1 port map( B1 => n1961_port, B2 => n11446, A => n11167, ZN 
                           => N2323);
   U15945 : OAI21_X1 port map( B1 => n1960_port, B2 => n11446, A => n11171, ZN 
                           => N2324);
   U15946 : OAI21_X1 port map( B1 => n1959_port, B2 => n11446, A => n11175, ZN 
                           => N2325);
   U15947 : OAI21_X1 port map( B1 => n1958_port, B2 => n11445, A => n11179, ZN 
                           => N2326);
   U15948 : OAI21_X1 port map( B1 => n1957_port, B2 => n11445, A => n11183, ZN 
                           => N2327);
   U15949 : OAI21_X1 port map( B1 => n1956_port, B2 => n11445, A => n11187, ZN 
                           => N2328);
   U15950 : OAI21_X1 port map( B1 => n1955_port, B2 => n11445, A => n11191, ZN 
                           => N2329);
   U15951 : OAI21_X1 port map( B1 => n1954_port, B2 => n11445, A => n11195, ZN 
                           => N2330);
   U15952 : OAI21_X1 port map( B1 => n1953_port, B2 => n11445, A => n11199, ZN 
                           => N2331);
   U15953 : OAI21_X1 port map( B1 => n1952_port, B2 => n11445, A => n11203, ZN 
                           => N2332);
   U15954 : OAI21_X1 port map( B1 => n1951_port, B2 => n11445, A => n11207, ZN 
                           => N2333);
   U15955 : OAI21_X1 port map( B1 => n1950_port, B2 => n11445, A => n11211, ZN 
                           => N2334);
   U15956 : OAI21_X1 port map( B1 => n1949_port, B2 => n11445, A => n11215, ZN 
                           => N2335);
   U15957 : OAI21_X1 port map( B1 => n1948_port, B2 => n11445, A => n11219, ZN 
                           => N2336);
   U15958 : OAI21_X1 port map( B1 => n1947_port, B2 => n11445, A => n11223, ZN 
                           => N2337);
   U15959 : OAI21_X1 port map( B1 => n1946_port, B2 => n11444, A => n11227, ZN 
                           => N2338);
   U15960 : OAI21_X1 port map( B1 => n1945_port, B2 => n11444, A => n11231, ZN 
                           => N2339);
   U15961 : OAI21_X1 port map( B1 => n1944_port, B2 => n11444, A => n11235, ZN 
                           => N2340);
   U15962 : OAI21_X1 port map( B1 => n1943_port, B2 => n11444, A => n11239, ZN 
                           => N2341);
   U15963 : OAI21_X1 port map( B1 => n1942_port, B2 => n11444, A => n11243, ZN 
                           => N2342);
   U15964 : OAI21_X1 port map( B1 => n1941_port, B2 => n11444, A => n11247, ZN 
                           => N2343);
   U15965 : OAI21_X1 port map( B1 => n1940_port, B2 => n11444, A => n11251, ZN 
                           => N2344);
   U15966 : OAI21_X1 port map( B1 => n1939_port, B2 => n11444, A => n11255, ZN 
                           => N2345);
   U15967 : OAI21_X1 port map( B1 => n1938_port, B2 => n11444, A => n11259, ZN 
                           => N2346);
   U15968 : OAI21_X1 port map( B1 => n1937_port, B2 => n11444, A => n11263, ZN 
                           => N2347);
   U15969 : OAI21_X1 port map( B1 => n1936_port, B2 => n11444, A => n11267, ZN 
                           => N2348);
   U15970 : OAI21_X1 port map( B1 => n1935_port, B2 => n11444, A => n11271, ZN 
                           => N2349);
   U15971 : OAI21_X1 port map( B1 => n1934_port, B2 => n11443, A => n11275, ZN 
                           => N2350);
   U15972 : OAI21_X1 port map( B1 => n1933_port, B2 => n11443, A => n11279, ZN 
                           => N2351);
   U15973 : OAI21_X1 port map( B1 => n1932_port, B2 => n11443, A => n11283, ZN 
                           => N2352);
   U15974 : OAI21_X1 port map( B1 => n1931_port, B2 => n11443, A => n11287, ZN 
                           => N2353);
   U15975 : OAI21_X1 port map( B1 => n1930_port, B2 => n11443, A => n11291, ZN 
                           => N2354);
   U15976 : OAI21_X1 port map( B1 => n1929_port, B2 => n11443, A => n11295, ZN 
                           => N2355);
   U15977 : OAI21_X1 port map( B1 => n1928_port, B2 => n11443, A => n11299, ZN 
                           => N2356);
   U15978 : OAI21_X1 port map( B1 => n1927_port, B2 => n11443, A => n11303, ZN 
                           => N2357);
   U15979 : OAI21_X1 port map( B1 => n1926_port, B2 => n11443, A => n11307, ZN 
                           => N2358);
   U15980 : OAI21_X1 port map( B1 => n1925_port, B2 => n11443, A => n11311, ZN 
                           => N2359);
   U15981 : OAI21_X1 port map( B1 => n1924_port, B2 => n11443, A => n11315, ZN 
                           => N2360);
   U15982 : OAI21_X1 port map( B1 => n1923_port, B2 => n11443, A => n11319, ZN 
                           => N2361);
   U15983 : OAI21_X1 port map( B1 => n1922_port, B2 => n11442, A => n11323, ZN 
                           => N2362);
   U15984 : OAI21_X1 port map( B1 => n1921_port, B2 => n11442, A => n11327, ZN 
                           => N2363);
   U15985 : OAI21_X1 port map( B1 => n1920_port, B2 => n11448, A => n11075, ZN 
                           => N2365);
   U15986 : OAI21_X1 port map( B1 => n1919_port, B2 => n11464, A => n11079, ZN 
                           => N2366);
   U15987 : OAI21_X1 port map( B1 => n1918_port, B2 => n11464, A => n11083, ZN 
                           => N2367);
   U15988 : OAI21_X1 port map( B1 => n1917_port, B2 => n11464, A => n11087, ZN 
                           => N2368);
   U15989 : OAI21_X1 port map( B1 => n1916_port, B2 => n11463, A => n11091, ZN 
                           => N2369);
   U15990 : OAI21_X1 port map( B1 => n1915_port, B2 => n11463, A => n11095, ZN 
                           => N2370);
   U15991 : OAI21_X1 port map( B1 => n1914_port, B2 => n11463, A => n11099, ZN 
                           => N2371);
   U15992 : OAI21_X1 port map( B1 => n1913_port, B2 => n11463, A => n11103, ZN 
                           => N2372);
   U15993 : OAI21_X1 port map( B1 => n1912_port, B2 => n11463, A => n11107, ZN 
                           => N2373);
   U15994 : OAI21_X1 port map( B1 => n1911_port, B2 => n11463, A => n11111, ZN 
                           => N2374);
   U15995 : OAI21_X1 port map( B1 => n1910_port, B2 => n11463, A => n11115, ZN 
                           => N2375);
   U15996 : OAI21_X1 port map( B1 => n1909_port, B2 => n11463, A => n11119, ZN 
                           => N2376);
   U15997 : OAI21_X1 port map( B1 => n1908_port, B2 => n11463, A => n11123, ZN 
                           => N2377);
   U15998 : OAI21_X1 port map( B1 => n1907_port, B2 => n11463, A => n11127, ZN 
                           => N2378);
   U15999 : OAI21_X1 port map( B1 => n1906_port, B2 => n11463, A => n11131, ZN 
                           => N2379);
   U16000 : OAI21_X1 port map( B1 => n1905_port, B2 => n11463, A => n11135, ZN 
                           => N2380);
   U16001 : OAI21_X1 port map( B1 => n1904_port, B2 => n11462, A => n11139, ZN 
                           => N2381);
   U16002 : OAI21_X1 port map( B1 => n1903_port, B2 => n11462, A => n11143, ZN 
                           => N2382);
   U16003 : OAI21_X1 port map( B1 => n1902_port, B2 => n11462, A => n11147, ZN 
                           => N2383);
   U16004 : OAI21_X1 port map( B1 => n1901_port, B2 => n11462, A => n11151, ZN 
                           => N2384);
   U16005 : OAI21_X1 port map( B1 => n1900_port, B2 => n11462, A => n11155, ZN 
                           => N2385);
   U16006 : OAI21_X1 port map( B1 => n1899_port, B2 => n11462, A => n11159, ZN 
                           => N2386);
   U16007 : OAI21_X1 port map( B1 => n1898_port, B2 => n11462, A => n11163, ZN 
                           => N2387);
   U16008 : OAI21_X1 port map( B1 => n1897_port, B2 => n11462, A => n11167, ZN 
                           => N2388);
   U16009 : OAI21_X1 port map( B1 => n1896_port, B2 => n11462, A => n11171, ZN 
                           => N2389);
   U16010 : OAI21_X1 port map( B1 => n1895_port, B2 => n11462, A => n11175, ZN 
                           => N2390);
   U16011 : OAI21_X1 port map( B1 => n1894_port, B2 => n11462, A => n11179, ZN 
                           => N2391);
   U16012 : OAI21_X1 port map( B1 => n1893_port, B2 => n11462, A => n11183, ZN 
                           => N2392);
   U16013 : OAI21_X1 port map( B1 => n1892_port, B2 => n11461, A => n11187, ZN 
                           => N2393);
   U16014 : OAI21_X1 port map( B1 => n1891_port, B2 => n11461, A => n11191, ZN 
                           => N2394);
   U16015 : OAI21_X1 port map( B1 => n1890_port, B2 => n11461, A => n11195, ZN 
                           => N2395);
   U16016 : OAI21_X1 port map( B1 => n1889_port, B2 => n11461, A => n11199, ZN 
                           => N2396);
   U16017 : OAI21_X1 port map( B1 => n1888_port, B2 => n11461, A => n11203, ZN 
                           => N2397);
   U16018 : OAI21_X1 port map( B1 => n1887_port, B2 => n11461, A => n11207, ZN 
                           => N2398);
   U16019 : OAI21_X1 port map( B1 => n1886_port, B2 => n11461, A => n11211, ZN 
                           => N2399);
   U16020 : OAI21_X1 port map( B1 => n1885_port, B2 => n11461, A => n11215, ZN 
                           => N2400);
   U16021 : OAI21_X1 port map( B1 => n1884_port, B2 => n11461, A => n11219, ZN 
                           => N2401);
   U16022 : OAI21_X1 port map( B1 => n1883_port, B2 => n11461, A => n11223, ZN 
                           => N2402);
   U16023 : OAI21_X1 port map( B1 => n1882_port, B2 => n11461, A => n11227, ZN 
                           => N2403);
   U16024 : OAI21_X1 port map( B1 => n1881_port, B2 => n11461, A => n11231, ZN 
                           => N2404);
   U16025 : OAI21_X1 port map( B1 => n1880_port, B2 => n11460, A => n11235, ZN 
                           => N2405);
   U16026 : OAI21_X1 port map( B1 => n1879_port, B2 => n11460, A => n11239, ZN 
                           => N2406);
   U16027 : OAI21_X1 port map( B1 => n1878_port, B2 => n11460, A => n11243, ZN 
                           => N2407);
   U16028 : OAI21_X1 port map( B1 => n1877_port, B2 => n11460, A => n11247, ZN 
                           => N2408);
   U16029 : OAI21_X1 port map( B1 => n1876_port, B2 => n11460, A => n11251, ZN 
                           => N2409);
   U16030 : OAI21_X1 port map( B1 => n1875_port, B2 => n11460, A => n11255, ZN 
                           => N2410);
   U16031 : OAI21_X1 port map( B1 => n1874_port, B2 => n11460, A => n11259, ZN 
                           => N2411);
   U16032 : OAI21_X1 port map( B1 => n1873_port, B2 => n11460, A => n11263, ZN 
                           => N2412);
   U16033 : OAI21_X1 port map( B1 => n1872_port, B2 => n11460, A => n11267, ZN 
                           => N2413);
   U16034 : OAI21_X1 port map( B1 => n1871_port, B2 => n11460, A => n11271, ZN 
                           => N2414);
   U16035 : OAI21_X1 port map( B1 => n1870_port, B2 => n11460, A => n11275, ZN 
                           => N2415);
   U16036 : OAI21_X1 port map( B1 => n1869_port, B2 => n11460, A => n11279, ZN 
                           => N2416);
   U16037 : OAI21_X1 port map( B1 => n1868_port, B2 => n11459, A => n11283, ZN 
                           => N2417);
   U16038 : OAI21_X1 port map( B1 => n1867_port, B2 => n11459, A => n11287, ZN 
                           => N2418);
   U16039 : OAI21_X1 port map( B1 => n1866_port, B2 => n11459, A => n11291, ZN 
                           => N2419);
   U16040 : OAI21_X1 port map( B1 => n1865_port, B2 => n11459, A => n11295, ZN 
                           => N2420);
   U16041 : OAI21_X1 port map( B1 => n1864_port, B2 => n11459, A => n11299, ZN 
                           => N2421);
   U16042 : OAI21_X1 port map( B1 => n1863_port, B2 => n11459, A => n11303, ZN 
                           => N2422);
   U16043 : OAI21_X1 port map( B1 => n1862_port, B2 => n11459, A => n11307, ZN 
                           => N2423);
   U16044 : OAI21_X1 port map( B1 => n1861_port, B2 => n11459, A => n11311, ZN 
                           => N2424);
   U16045 : OAI21_X1 port map( B1 => n1860_port, B2 => n11459, A => n11315, ZN 
                           => N2425);
   U16046 : OAI21_X1 port map( B1 => n1859_port, B2 => n11459, A => n11319, ZN 
                           => N2426);
   U16047 : OAI21_X1 port map( B1 => n1858_port, B2 => n11459, A => n11323, ZN 
                           => N2427);
   U16048 : OAI21_X1 port map( B1 => n1857_port, B2 => n11459, A => n11327, ZN 
                           => N2428);
   U16049 : OAI21_X1 port map( B1 => n1856_port, B2 => n11458, A => n11075, ZN 
                           => N2430);
   U16050 : OAI21_X1 port map( B1 => n1855_port, B2 => n11458, A => n11079, ZN 
                           => N2431);
   U16051 : OAI21_X1 port map( B1 => n1854_port, B2 => n11458, A => n11083, ZN 
                           => N2432);
   U16052 : OAI21_X1 port map( B1 => n1853_port, B2 => n11458, A => n11087, ZN 
                           => N2433);
   U16053 : OAI21_X1 port map( B1 => n1852_port, B2 => n11458, A => n11091, ZN 
                           => N2434);
   U16054 : OAI21_X1 port map( B1 => n1851_port, B2 => n11458, A => n11095, ZN 
                           => N2435);
   U16055 : OAI21_X1 port map( B1 => n1850_port, B2 => n11458, A => n11099, ZN 
                           => N2436);
   U16056 : OAI21_X1 port map( B1 => n1849_port, B2 => n11458, A => n11103, ZN 
                           => N2437);
   U16057 : OAI21_X1 port map( B1 => n1848_port, B2 => n11458, A => n11107, ZN 
                           => N2438);
   U16058 : OAI21_X1 port map( B1 => n1847_port, B2 => n11458, A => n11111, ZN 
                           => N2439);
   U16059 : OAI21_X1 port map( B1 => n1846_port, B2 => n11458, A => n11115, ZN 
                           => N2440);
   U16060 : OAI21_X1 port map( B1 => n1845_port, B2 => n11457, A => n11119, ZN 
                           => N2441);
   U16061 : OAI21_X1 port map( B1 => n1844_port, B2 => n11457, A => n11123, ZN 
                           => N2442);
   U16062 : OAI21_X1 port map( B1 => n1843_port, B2 => n11457, A => n11127, ZN 
                           => N2443);
   U16063 : OAI21_X1 port map( B1 => n1842_port, B2 => n11457, A => n11131, ZN 
                           => N2444);
   U16064 : OAI21_X1 port map( B1 => n1841_port, B2 => n11457, A => n11135, ZN 
                           => N2445);
   U16065 : OAI21_X1 port map( B1 => n1840_port, B2 => n11457, A => n11139, ZN 
                           => N2446);
   U16066 : OAI21_X1 port map( B1 => n1839_port, B2 => n11457, A => n11143, ZN 
                           => N2447);
   U16067 : OAI21_X1 port map( B1 => n1838_port, B2 => n11457, A => n11147, ZN 
                           => N2448);
   U16068 : OAI21_X1 port map( B1 => n1837_port, B2 => n11457, A => n11151, ZN 
                           => N2449);
   U16069 : OAI21_X1 port map( B1 => n1836_port, B2 => n11457, A => n11155, ZN 
                           => N2450);
   U16070 : OAI21_X1 port map( B1 => n1835_port, B2 => n11457, A => n11159, ZN 
                           => N2451);
   U16071 : OAI21_X1 port map( B1 => n1834_port, B2 => n11457, A => n11163, ZN 
                           => N2452);
   U16072 : OAI21_X1 port map( B1 => n1833_port, B2 => n11456, A => n11167, ZN 
                           => N2453);
   U16073 : OAI21_X1 port map( B1 => n1832_port, B2 => n11456, A => n11171, ZN 
                           => N2454);
   U16074 : OAI21_X1 port map( B1 => n1831_port, B2 => n11456, A => n11175, ZN 
                           => N2455);
   U16075 : OAI21_X1 port map( B1 => n1830_port, B2 => n11456, A => n11179, ZN 
                           => N2456);
   U16076 : OAI21_X1 port map( B1 => n1829_port, B2 => n11456, A => n11183, ZN 
                           => N2457);
   U16077 : OAI21_X1 port map( B1 => n1828_port, B2 => n11456, A => n11187, ZN 
                           => N2458);
   U16078 : OAI21_X1 port map( B1 => n1827_port, B2 => n11456, A => n11191, ZN 
                           => N2459);
   U16079 : OAI21_X1 port map( B1 => n1826_port, B2 => n11456, A => n11195, ZN 
                           => N2460);
   U16080 : OAI21_X1 port map( B1 => n1825_port, B2 => n11456, A => n11199, ZN 
                           => N2461);
   U16081 : OAI21_X1 port map( B1 => n1824_port, B2 => n11456, A => n11203, ZN 
                           => N2462);
   U16082 : OAI21_X1 port map( B1 => n1823_port, B2 => n11456, A => n11207, ZN 
                           => N2463);
   U16083 : OAI21_X1 port map( B1 => n1822_port, B2 => n11456, A => n11211, ZN 
                           => N2464);
   U16084 : OAI21_X1 port map( B1 => n1821_port, B2 => n11455, A => n11215, ZN 
                           => N2465);
   U16085 : OAI21_X1 port map( B1 => n1820_port, B2 => n11455, A => n11219, ZN 
                           => N2466);
   U16086 : OAI21_X1 port map( B1 => n1819_port, B2 => n11455, A => n11223, ZN 
                           => N2467);
   U16087 : OAI21_X1 port map( B1 => n1818_port, B2 => n11455, A => n11227, ZN 
                           => N2468);
   U16088 : OAI21_X1 port map( B1 => n1817_port, B2 => n11455, A => n11231, ZN 
                           => N2469);
   U16089 : OAI21_X1 port map( B1 => n1816_port, B2 => n11455, A => n11235, ZN 
                           => N2470);
   U16090 : OAI21_X1 port map( B1 => n1815_port, B2 => n11455, A => n11239, ZN 
                           => N2471);
   U16091 : OAI21_X1 port map( B1 => n1814_port, B2 => n11455, A => n11243, ZN 
                           => N2472);
   U16092 : OAI21_X1 port map( B1 => n1813_port, B2 => n11455, A => n11247, ZN 
                           => N2473);
   U16093 : OAI21_X1 port map( B1 => n1812_port, B2 => n11455, A => n11251, ZN 
                           => N2474);
   U16094 : OAI21_X1 port map( B1 => n1811_port, B2 => n11455, A => n11255, ZN 
                           => N2475);
   U16095 : OAI21_X1 port map( B1 => n1810_port, B2 => n11455, A => n11259, ZN 
                           => N2476);
   U16096 : OAI21_X1 port map( B1 => n1809_port, B2 => n11454, A => n11263, ZN 
                           => N2477);
   U16097 : OAI21_X1 port map( B1 => n1808_port, B2 => n11454, A => n11267, ZN 
                           => N2478);
   U16098 : OAI21_X1 port map( B1 => n1807_port, B2 => n11454, A => n11271, ZN 
                           => N2479);
   U16099 : OAI21_X1 port map( B1 => n1806_port, B2 => n11454, A => n11275, ZN 
                           => N2480);
   U16100 : OAI21_X1 port map( B1 => n1805_port, B2 => n11454, A => n11279, ZN 
                           => N2481);
   U16101 : OAI21_X1 port map( B1 => n1804_port, B2 => n11454, A => n11283, ZN 
                           => N2482);
   U16102 : OAI21_X1 port map( B1 => n1803_port, B2 => n11454, A => n11287, ZN 
                           => N2483);
   U16103 : OAI21_X1 port map( B1 => n1802_port, B2 => n11454, A => n11291, ZN 
                           => N2484);
   U16104 : OAI21_X1 port map( B1 => n1801_port, B2 => n11454, A => n11295, ZN 
                           => N2485);
   U16105 : OAI21_X1 port map( B1 => n1800_port, B2 => n11454, A => n11299, ZN 
                           => N2486);
   U16106 : OAI21_X1 port map( B1 => n1799_port, B2 => n11454, A => n11303, ZN 
                           => N2487);
   U16107 : OAI21_X1 port map( B1 => n1798_port, B2 => n11454, A => n11307, ZN 
                           => N2488);
   U16108 : OAI21_X1 port map( B1 => n1797_port, B2 => n11453, A => n11311, ZN 
                           => N2489);
   U16109 : OAI21_X1 port map( B1 => n1796_port, B2 => n11453, A => n11315, ZN 
                           => N2490);
   U16110 : OAI21_X1 port map( B1 => n1795_port, B2 => n11453, A => n11319, ZN 
                           => N2491);
   U16111 : OAI21_X1 port map( B1 => n1794_port, B2 => n11464, A => n11323, ZN 
                           => N2492);
   U16112 : OAI21_X1 port map( B1 => n1793_port, B2 => n11453, A => n11327, ZN 
                           => N2493);
   U16113 : OAI21_X1 port map( B1 => n1792_port, B2 => n11453, A => n11075, ZN 
                           => N2495);
   U16114 : OAI21_X1 port map( B1 => n1791_port, B2 => n11458, A => n11079, ZN 
                           => N2496);
   U16115 : OAI21_X1 port map( B1 => n1790_port, B2 => n11432, A => n11083, ZN 
                           => N2497);
   U16116 : OAI21_X1 port map( B1 => n1789_port, B2 => n11431, A => n11087, ZN 
                           => N2498);
   U16117 : OAI21_X1 port map( B1 => n1788_port, B2 => n11431, A => n11091, ZN 
                           => N2499);
   U16118 : OAI21_X1 port map( B1 => n1787_port, B2 => n11431, A => n11095, ZN 
                           => N2500);
   U16119 : OAI21_X1 port map( B1 => n1786_port, B2 => n11431, A => n11099, ZN 
                           => N2501);
   U16120 : OAI21_X1 port map( B1 => n1785_port, B2 => n11431, A => n11103, ZN 
                           => N2502);
   U16121 : OAI21_X1 port map( B1 => n1784_port, B2 => n11431, A => n11107, ZN 
                           => N2503);
   U16122 : OAI21_X1 port map( B1 => n1783_port, B2 => n11431, A => n11111, ZN 
                           => N2504);
   U16123 : OAI21_X1 port map( B1 => n1782_port, B2 => n11431, A => n11115, ZN 
                           => N2505);
   U16124 : OAI21_X1 port map( B1 => n1781_port, B2 => n11431, A => n11119, ZN 
                           => N2506);
   U16125 : OAI21_X1 port map( B1 => n1780_port, B2 => n11431, A => n11123, ZN 
                           => N2507);
   U16126 : OAI21_X1 port map( B1 => n1779_port, B2 => n11431, A => n11127, ZN 
                           => N2508);
   U16127 : OAI21_X1 port map( B1 => n1778_port, B2 => n11431, A => n11131, ZN 
                           => N2509);
   U16128 : OAI21_X1 port map( B1 => n1777_port, B2 => n11430, A => n11135, ZN 
                           => N2510);
   U16129 : OAI21_X1 port map( B1 => n1776_port, B2 => n11430, A => n11139, ZN 
                           => N2511);
   U16130 : OAI21_X1 port map( B1 => n1775_port, B2 => n11430, A => n11143, ZN 
                           => N2512);
   U16131 : OAI21_X1 port map( B1 => n1774_port, B2 => n11430, A => n11147, ZN 
                           => N2513);
   U16132 : OAI21_X1 port map( B1 => n1773_port, B2 => n11430, A => n11151, ZN 
                           => N2514);
   U16133 : OAI21_X1 port map( B1 => n1772_port, B2 => n11430, A => n11155, ZN 
                           => N2515);
   U16134 : OAI21_X1 port map( B1 => n1771_port, B2 => n11430, A => n11159, ZN 
                           => N2516);
   U16135 : OAI21_X1 port map( B1 => n1770_port, B2 => n11430, A => n11163, ZN 
                           => N2517);
   U16136 : OAI21_X1 port map( B1 => n1769_port, B2 => n11430, A => n11167, ZN 
                           => N2518);
   U16137 : OAI21_X1 port map( B1 => n1768_port, B2 => n11430, A => n11171, ZN 
                           => N2519);
   U16138 : OAI21_X1 port map( B1 => n1767_port, B2 => n11430, A => n11175, ZN 
                           => N2520);
   U16139 : OAI21_X1 port map( B1 => n1766_port, B2 => n11430, A => n11179, ZN 
                           => N2521);
   U16140 : OAI21_X1 port map( B1 => n1765_port, B2 => n11429, A => n11183, ZN 
                           => N2522);
   U16141 : OAI21_X1 port map( B1 => n1764_port, B2 => n11429, A => n11187, ZN 
                           => N2523);
   U16142 : OAI21_X1 port map( B1 => n1763_port, B2 => n11429, A => n11191, ZN 
                           => N2524);
   U16143 : OAI21_X1 port map( B1 => n1762_port, B2 => n11429, A => n11195, ZN 
                           => N2525);
   U16144 : OAI21_X1 port map( B1 => n1761_port, B2 => n11429, A => n11199, ZN 
                           => N2526);
   U16145 : OAI21_X1 port map( B1 => n1760_port, B2 => n11429, A => n11203, ZN 
                           => N2527);
   U16146 : OAI21_X1 port map( B1 => n1759_port, B2 => n11429, A => n11207, ZN 
                           => N2528);
   U16147 : OAI21_X1 port map( B1 => n1758_port, B2 => n11429, A => n11211, ZN 
                           => N2529);
   U16148 : OAI21_X1 port map( B1 => n1757_port, B2 => n11429, A => n11215, ZN 
                           => N2530);
   U16149 : OAI21_X1 port map( B1 => n1756_port, B2 => n11429, A => n11219, ZN 
                           => N2531);
   U16150 : OAI21_X1 port map( B1 => n1755_port, B2 => n11429, A => n11223, ZN 
                           => N2532);
   U16151 : OAI21_X1 port map( B1 => n1754_port, B2 => n11429, A => n11227, ZN 
                           => N2533);
   U16152 : OAI21_X1 port map( B1 => n1753_port, B2 => n11428, A => n11231, ZN 
                           => N2534);
   U16153 : OAI21_X1 port map( B1 => n1752_port, B2 => n11428, A => n11235, ZN 
                           => N2535);
   U16154 : OAI21_X1 port map( B1 => n1751_port, B2 => n11428, A => n11239, ZN 
                           => N2536);
   U16155 : OAI21_X1 port map( B1 => n1750_port, B2 => n11428, A => n11243, ZN 
                           => N2537);
   U16156 : OAI21_X1 port map( B1 => n1749_port, B2 => n11428, A => n11247, ZN 
                           => N2538);
   U16157 : OAI21_X1 port map( B1 => n1748_port, B2 => n11428, A => n11251, ZN 
                           => N2539);
   U16158 : OAI21_X1 port map( B1 => n1747_port, B2 => n11428, A => n11255, ZN 
                           => N2540);
   U16159 : OAI21_X1 port map( B1 => n1746_port, B2 => n11428, A => n11259, ZN 
                           => N2541);
   U16160 : OAI21_X1 port map( B1 => n1745_port, B2 => n11428, A => n11263, ZN 
                           => N2542);
   U16161 : OAI21_X1 port map( B1 => n1744_port, B2 => n11428, A => n11267, ZN 
                           => N2543);
   U16162 : OAI21_X1 port map( B1 => n1743_port, B2 => n11428, A => n11271, ZN 
                           => N2544);
   U16163 : OAI21_X1 port map( B1 => n1742_port, B2 => n11428, A => n11275, ZN 
                           => N2545);
   U16164 : OAI21_X1 port map( B1 => n1741_port, B2 => n11427, A => n11279, ZN 
                           => N2546);
   U16165 : OAI21_X1 port map( B1 => n1740_port, B2 => n11427, A => n11283, ZN 
                           => N2547);
   U16166 : OAI21_X1 port map( B1 => n1739_port, B2 => n11427, A => n11287, ZN 
                           => N2548);
   U16167 : OAI21_X1 port map( B1 => n1738_port, B2 => n11427, A => n11291, ZN 
                           => N2549);
   U16168 : OAI21_X1 port map( B1 => n1737_port, B2 => n11427, A => n11295, ZN 
                           => N2550);
   U16169 : OAI21_X1 port map( B1 => n1736_port, B2 => n11427, A => n11299, ZN 
                           => N2551);
   U16170 : OAI21_X1 port map( B1 => n1735_port, B2 => n11427, A => n11303, ZN 
                           => N2552);
   U16171 : OAI21_X1 port map( B1 => n1734_port, B2 => n11427, A => n11307, ZN 
                           => N2553);
   U16172 : OAI21_X1 port map( B1 => n1733_port, B2 => n11427, A => n11311, ZN 
                           => N2554);
   U16173 : OAI21_X1 port map( B1 => n1732_port, B2 => n11427, A => n11315, ZN 
                           => N2555);
   U16174 : OAI21_X1 port map( B1 => n1731_port, B2 => n11427, A => n11319, ZN 
                           => N2556);
   U16175 : OAI21_X1 port map( B1 => n1730_port, B2 => n11427, A => n11323, ZN 
                           => N2557);
   U16176 : OAI21_X1 port map( B1 => n1729_port, B2 => n11426, A => n11327, ZN 
                           => N2558);
   U16177 : OAI21_X1 port map( B1 => n1728_port, B2 => n11426, A => n11075, ZN 
                           => N2560);
   U16178 : OAI21_X1 port map( B1 => n1727_port, B2 => n11426, A => n11079, ZN 
                           => N2561);
   U16179 : OAI21_X1 port map( B1 => n1726_port, B2 => n11426, A => n11083, ZN 
                           => N2562);
   U16180 : OAI21_X1 port map( B1 => n1725_port, B2 => n11426, A => n11087, ZN 
                           => N2563);
   U16181 : OAI21_X1 port map( B1 => n1724_port, B2 => n11426, A => n11091, ZN 
                           => N2564);
   U16182 : OAI21_X1 port map( B1 => n1723_port, B2 => n11426, A => n11095, ZN 
                           => N2565);
   U16183 : OAI21_X1 port map( B1 => n1722_port, B2 => n11426, A => n11099, ZN 
                           => N2566);
   U16184 : OAI21_X1 port map( B1 => n1721_port, B2 => n11426, A => n11103, ZN 
                           => N2567);
   U16185 : OAI21_X1 port map( B1 => n1720_port, B2 => n11426, A => n11107, ZN 
                           => N2568);
   U16186 : OAI21_X1 port map( B1 => n1719_port, B2 => n11426, A => n11111, ZN 
                           => N2569);
   U16187 : OAI21_X1 port map( B1 => n1718_port, B2 => n11425, A => n11115, ZN 
                           => N2570);
   U16188 : OAI21_X1 port map( B1 => n1717_port, B2 => n11425, A => n11119, ZN 
                           => N2571);
   U16189 : OAI21_X1 port map( B1 => n1716_port, B2 => n11425, A => n11123, ZN 
                           => N2572);
   U16190 : OAI21_X1 port map( B1 => n1715_port, B2 => n11425, A => n11127, ZN 
                           => N2573);
   U16191 : OAI21_X1 port map( B1 => n1714_port, B2 => n11425, A => n11131, ZN 
                           => N2574);
   U16192 : OAI21_X1 port map( B1 => n1713_port, B2 => n11425, A => n11135, ZN 
                           => N2575);
   U16193 : OAI21_X1 port map( B1 => n1712_port, B2 => n11425, A => n11139, ZN 
                           => N2576);
   U16194 : OAI21_X1 port map( B1 => n1711_port, B2 => n11425, A => n11143, ZN 
                           => N2577);
   U16195 : OAI21_X1 port map( B1 => n1710_port, B2 => n11425, A => n11147, ZN 
                           => N2578);
   U16196 : OAI21_X1 port map( B1 => n1709_port, B2 => n11425, A => n11151, ZN 
                           => N2579);
   U16197 : OAI21_X1 port map( B1 => n1708_port, B2 => n11425, A => n11155, ZN 
                           => N2580);
   U16198 : OAI21_X1 port map( B1 => n1707_port, B2 => n11425, A => n11159, ZN 
                           => N2581);
   U16199 : OAI21_X1 port map( B1 => n1706_port, B2 => n11424, A => n11163, ZN 
                           => N2582);
   U16200 : OAI21_X1 port map( B1 => n1705_port, B2 => n11424, A => n11167, ZN 
                           => N2583);
   U16201 : OAI21_X1 port map( B1 => n1704_port, B2 => n11424, A => n11171, ZN 
                           => N2584);
   U16202 : OAI21_X1 port map( B1 => n1703_port, B2 => n11424, A => n11175, ZN 
                           => N2585);
   U16203 : OAI21_X1 port map( B1 => n1702_port, B2 => n11424, A => n11179, ZN 
                           => N2586);
   U16204 : OAI21_X1 port map( B1 => n1701_port, B2 => n11424, A => n11183, ZN 
                           => N2587);
   U16205 : OAI21_X1 port map( B1 => n1700_port, B2 => n11424, A => n11187, ZN 
                           => N2588);
   U16206 : OAI21_X1 port map( B1 => n1699_port, B2 => n11424, A => n11191, ZN 
                           => N2589);
   U16207 : OAI21_X1 port map( B1 => n1698_port, B2 => n11424, A => n11195, ZN 
                           => N2590);
   U16208 : OAI21_X1 port map( B1 => n1697_port, B2 => n11424, A => n11199, ZN 
                           => N2591);
   U16209 : OAI21_X1 port map( B1 => n1696_port, B2 => n11424, A => n11203, ZN 
                           => N2592);
   U16210 : OAI21_X1 port map( B1 => n1695_port, B2 => n11424, A => n11207, ZN 
                           => N2593);
   U16211 : OAI21_X1 port map( B1 => n1694_port, B2 => n11423, A => n11211, ZN 
                           => N2594);
   U16212 : OAI21_X1 port map( B1 => n1693_port, B2 => n11423, A => n11215, ZN 
                           => N2595);
   U16213 : OAI21_X1 port map( B1 => n1692_port, B2 => n11423, A => n11219, ZN 
                           => N2596);
   U16214 : OAI21_X1 port map( B1 => n1691_port, B2 => n11423, A => n11223, ZN 
                           => N2597);
   U16215 : OAI21_X1 port map( B1 => n1690_port, B2 => n11423, A => n11227, ZN 
                           => N2598);
   U16216 : OAI21_X1 port map( B1 => n1689_port, B2 => n11423, A => n11231, ZN 
                           => N2599);
   U16217 : OAI21_X1 port map( B1 => n1688_port, B2 => n11423, A => n11235, ZN 
                           => N2600);
   U16218 : OAI21_X1 port map( B1 => n1687_port, B2 => n11423, A => n11239, ZN 
                           => N2601);
   U16219 : OAI21_X1 port map( B1 => n1686_port, B2 => n11423, A => n11243, ZN 
                           => N2602);
   U16220 : OAI21_X1 port map( B1 => n1685_port, B2 => n11423, A => n11247, ZN 
                           => N2603);
   U16221 : OAI21_X1 port map( B1 => n1684_port, B2 => n11423, A => n11251, ZN 
                           => N2604);
   U16222 : OAI21_X1 port map( B1 => n1683_port, B2 => n11423, A => n11255, ZN 
                           => N2605);
   U16223 : OAI21_X1 port map( B1 => n1682_port, B2 => n11422, A => n11259, ZN 
                           => N2606);
   U16224 : OAI21_X1 port map( B1 => n1681_port, B2 => n11422, A => n11263, ZN 
                           => N2607);
   U16225 : OAI21_X1 port map( B1 => n1680_port, B2 => n11422, A => n11267, ZN 
                           => N2608);
   U16226 : OAI21_X1 port map( B1 => n1679_port, B2 => n11422, A => n11271, ZN 
                           => N2609);
   U16227 : OAI21_X1 port map( B1 => n1678_port, B2 => n11422, A => n11275, ZN 
                           => N2610);
   U16228 : OAI21_X1 port map( B1 => n1677_port, B2 => n11422, A => n11279, ZN 
                           => N2611);
   U16229 : OAI21_X1 port map( B1 => n1676_port, B2 => n11422, A => n11283, ZN 
                           => N2612);
   U16230 : OAI21_X1 port map( B1 => n1675_port, B2 => n11422, A => n11287, ZN 
                           => N2613);
   U16231 : OAI21_X1 port map( B1 => n1674_port, B2 => n11422, A => n11291, ZN 
                           => N2614);
   U16232 : OAI21_X1 port map( B1 => n1673_port, B2 => n11422, A => n11295, ZN 
                           => N2615);
   U16233 : OAI21_X1 port map( B1 => n1672_port, B2 => n11422, A => n11299, ZN 
                           => N2616);
   U16234 : OAI21_X1 port map( B1 => n1671_port, B2 => n11422, A => n11303, ZN 
                           => N2617);
   U16235 : OAI21_X1 port map( B1 => n1670_port, B2 => n11421, A => n11307, ZN 
                           => N2618);
   U16236 : OAI21_X1 port map( B1 => n1669_port, B2 => n11421, A => n11311, ZN 
                           => N2619);
   U16237 : OAI21_X1 port map( B1 => n1668_port, B2 => n11421, A => n11315, ZN 
                           => N2620);
   U16238 : OAI21_X1 port map( B1 => n1667_port, B2 => n11421, A => n11319, ZN 
                           => N2621);
   U16239 : OAI21_X1 port map( B1 => n1666_port, B2 => n11421, A => n11323, ZN 
                           => N2622);
   U16240 : OAI21_X1 port map( B1 => n1665_port, B2 => n11421, A => n11327, ZN 
                           => N2623);
   U16241 : OAI21_X1 port map( B1 => n1664_port, B2 => n11421, A => n11075, ZN 
                           => N2625);
   U16242 : OAI21_X1 port map( B1 => n1663_port, B2 => n11421, A => n11079, ZN 
                           => N2626);
   U16243 : OAI21_X1 port map( B1 => n1662_port, B2 => n11426, A => n11083, ZN 
                           => N2627);
   U16244 : OAI21_X1 port map( B1 => n1661_port, B2 => n11442, A => n11087, ZN 
                           => N2628);
   U16245 : OAI21_X1 port map( B1 => n1660_port, B2 => n11442, A => n11091, ZN 
                           => N2629);
   U16246 : OAI21_X1 port map( B1 => n1659_port, B2 => n11442, A => n11095, ZN 
                           => N2630);
   U16247 : OAI21_X1 port map( B1 => n1658_port, B2 => n11442, A => n11099, ZN 
                           => N2631);
   U16248 : OAI21_X1 port map( B1 => n1657_port, B2 => n11442, A => n11103, ZN 
                           => N2632);
   U16249 : OAI21_X1 port map( B1 => n1656_port, B2 => n11442, A => n11107, ZN 
                           => N2633);
   U16250 : OAI21_X1 port map( B1 => n1655_port, B2 => n11442, A => n11111, ZN 
                           => N2634);
   U16251 : OAI21_X1 port map( B1 => n1654_port, B2 => n11442, A => n11115, ZN 
                           => N2635);
   U16252 : OAI21_X1 port map( B1 => n1653_port, B2 => n11442, A => n11119, ZN 
                           => N2636);
   U16253 : OAI21_X1 port map( B1 => n1652_port, B2 => n11441, A => n11123, ZN 
                           => N2637);
   U16254 : OAI21_X1 port map( B1 => n1651_port, B2 => n11441, A => n11127, ZN 
                           => N2638);
   U16255 : OAI21_X1 port map( B1 => n1650_port, B2 => n11441, A => n11131, ZN 
                           => N2639);
   U16256 : OAI21_X1 port map( B1 => n1649_port, B2 => n11441, A => n11135, ZN 
                           => N2640);
   U16257 : OAI21_X1 port map( B1 => n1648_port, B2 => n11441, A => n11139, ZN 
                           => N2641);
   U16258 : OAI21_X1 port map( B1 => n1647_port, B2 => n11441, A => n11143, ZN 
                           => N2642);
   U16259 : OAI21_X1 port map( B1 => n1646_port, B2 => n11441, A => n11147, ZN 
                           => N2643);
   U16260 : OAI21_X1 port map( B1 => n1645_port, B2 => n11441, A => n11151, ZN 
                           => N2644);
   U16261 : OAI21_X1 port map( B1 => n1644_port, B2 => n11441, A => n11155, ZN 
                           => N2645);
   U16262 : OAI21_X1 port map( B1 => n1643_port, B2 => n11441, A => n11159, ZN 
                           => N2646);
   U16263 : OAI21_X1 port map( B1 => n1642_port, B2 => n11441, A => n11163, ZN 
                           => N2647);
   U16264 : OAI21_X1 port map( B1 => n1641_port, B2 => n11441, A => n11167, ZN 
                           => N2648);
   U16265 : OAI21_X1 port map( B1 => n1640_port, B2 => n11440, A => n11171, ZN 
                           => N2649);
   U16266 : OAI21_X1 port map( B1 => n1639_port, B2 => n11440, A => n11175, ZN 
                           => N2650);
   U16267 : OAI21_X1 port map( B1 => n1638_port, B2 => n11440, A => n11179, ZN 
                           => N2651);
   U16268 : OAI21_X1 port map( B1 => n1637_port, B2 => n11440, A => n11183, ZN 
                           => N2652);
   U16269 : OAI21_X1 port map( B1 => n1636_port, B2 => n11440, A => n11187, ZN 
                           => N2653);
   U16270 : OAI21_X1 port map( B1 => n1635_port, B2 => n11440, A => n11191, ZN 
                           => N2654);
   U16271 : OAI21_X1 port map( B1 => n1634_port, B2 => n11440, A => n11195, ZN 
                           => N2655);
   U16272 : OAI21_X1 port map( B1 => n1633_port, B2 => n11440, A => n11199, ZN 
                           => N2656);
   U16273 : OAI21_X1 port map( B1 => n1632_port, B2 => n11440, A => n11203, ZN 
                           => N2657);
   U16274 : OAI21_X1 port map( B1 => n1631_port, B2 => n11440, A => n11207, ZN 
                           => N2658);
   U16275 : OAI21_X1 port map( B1 => n1630_port, B2 => n11440, A => n11211, ZN 
                           => N2659);
   U16276 : OAI21_X1 port map( B1 => n1629_port, B2 => n11440, A => n11215, ZN 
                           => N2660);
   U16277 : OAI21_X1 port map( B1 => n1628_port, B2 => n11439, A => n11219, ZN 
                           => N2661);
   U16278 : OAI21_X1 port map( B1 => n1627_port, B2 => n11439, A => n11223, ZN 
                           => N2662);
   U16279 : OAI21_X1 port map( B1 => n1626_port, B2 => n11439, A => n11227, ZN 
                           => N2663);
   U16280 : OAI21_X1 port map( B1 => n1625_port, B2 => n11439, A => n11231, ZN 
                           => N2664);
   U16281 : OAI21_X1 port map( B1 => n1624_port, B2 => n11439, A => n11235, ZN 
                           => N2665);
   U16282 : OAI21_X1 port map( B1 => n1623_port, B2 => n11439, A => n11239, ZN 
                           => N2666);
   U16283 : OAI21_X1 port map( B1 => n1622_port, B2 => n11439, A => n11243, ZN 
                           => N2667);
   U16284 : OAI21_X1 port map( B1 => n1621_port, B2 => n11439, A => n11247, ZN 
                           => N2668);
   U16285 : OAI21_X1 port map( B1 => n1620_port, B2 => n11439, A => n11251, ZN 
                           => N2669);
   U16286 : OAI21_X1 port map( B1 => n1619_port, B2 => n11439, A => n11255, ZN 
                           => N2670);
   U16287 : OAI21_X1 port map( B1 => n1618_port, B2 => n11439, A => n11259, ZN 
                           => N2671);
   U16288 : OAI21_X1 port map( B1 => n1617_port, B2 => n11439, A => n11263, ZN 
                           => N2672);
   U16289 : OAI21_X1 port map( B1 => n1616_port, B2 => n11438, A => n11267, ZN 
                           => N2673);
   U16290 : OAI21_X1 port map( B1 => n1615_port, B2 => n11438, A => n11271, ZN 
                           => N2674);
   U16291 : OAI21_X1 port map( B1 => n1614_port, B2 => n11438, A => n11275, ZN 
                           => N2675);
   U16292 : OAI21_X1 port map( B1 => n1613_port, B2 => n11438, A => n11279, ZN 
                           => N2676);
   U16293 : OAI21_X1 port map( B1 => n1612_port, B2 => n11438, A => n11283, ZN 
                           => N2677);
   U16294 : OAI21_X1 port map( B1 => n1611_port, B2 => n11438, A => n11287, ZN 
                           => N2678);
   U16295 : OAI21_X1 port map( B1 => n1610_port, B2 => n11438, A => n11291, ZN 
                           => N2679);
   U16296 : OAI21_X1 port map( B1 => n1609_port, B2 => n11438, A => n11295, ZN 
                           => N2680);
   U16297 : OAI21_X1 port map( B1 => n1608_port, B2 => n11438, A => n11299, ZN 
                           => N2681);
   U16298 : OAI21_X1 port map( B1 => n1607_port, B2 => n11438, A => n11303, ZN 
                           => N2682);
   U16299 : OAI21_X1 port map( B1 => n1606_port, B2 => n11438, A => n11307, ZN 
                           => N2683);
   U16300 : OAI21_X1 port map( B1 => n1605_port, B2 => n11438, A => n11311, ZN 
                           => N2684);
   U16301 : OAI21_X1 port map( B1 => n1604_port, B2 => n11437, A => n11315, ZN 
                           => N2685);
   U16302 : OAI21_X1 port map( B1 => n1603_port, B2 => n11437, A => n11319, ZN 
                           => N2686);
   U16303 : OAI21_X1 port map( B1 => n1602_port, B2 => n11437, A => n11323, ZN 
                           => N2687);
   U16304 : OAI21_X1 port map( B1 => n1601_port, B2 => n11437, A => n11327, ZN 
                           => N2688);
   U16305 : OAI21_X1 port map( B1 => n1600_port, B2 => n11437, A => n11075, ZN 
                           => N2690);
   U16306 : OAI21_X1 port map( B1 => n1599_port, B2 => n11437, A => n11079, ZN 
                           => N2691);
   U16307 : OAI21_X1 port map( B1 => n1598_port, B2 => n11437, A => n11083, ZN 
                           => N2692);
   U16308 : OAI21_X1 port map( B1 => n1597_port, B2 => n11437, A => n11087, ZN 
                           => N2693);
   U16309 : OAI21_X1 port map( B1 => n1596_port, B2 => n11437, A => n11091, ZN 
                           => N2694);
   U16310 : OAI21_X1 port map( B1 => n1595_port, B2 => n11437, A => n11095, ZN 
                           => N2695);
   U16311 : OAI21_X1 port map( B1 => n1594_port, B2 => n11437, A => n11099, ZN 
                           => N2696);
   U16312 : OAI21_X1 port map( B1 => n1593_port, B2 => n11436, A => n11103, ZN 
                           => N2697);
   U16313 : OAI21_X1 port map( B1 => n1592_port, B2 => n11436, A => n11107, ZN 
                           => N2698);
   U16314 : OAI21_X1 port map( B1 => n1591_port, B2 => n11436, A => n11111, ZN 
                           => N2699);
   U16315 : OAI21_X1 port map( B1 => n1590_port, B2 => n11436, A => n11115, ZN 
                           => N2700);
   U16316 : OAI21_X1 port map( B1 => n1589_port, B2 => n11436, A => n11119, ZN 
                           => N2701);
   U16317 : OAI21_X1 port map( B1 => n1588_port, B2 => n11436, A => n11123, ZN 
                           => N2702);
   U16318 : OAI21_X1 port map( B1 => n1587_port, B2 => n11436, A => n11127, ZN 
                           => N2703);
   U16319 : OAI21_X1 port map( B1 => n1586_port, B2 => n11436, A => n11131, ZN 
                           => N2704);
   U16320 : OAI21_X1 port map( B1 => n1585_port, B2 => n11436, A => n11135, ZN 
                           => N2705);
   U16321 : OAI21_X1 port map( B1 => n1584_port, B2 => n11436, A => n11139, ZN 
                           => N2706);
   U16322 : OAI21_X1 port map( B1 => n1583_port, B2 => n11436, A => n11143, ZN 
                           => N2707);
   U16323 : OAI21_X1 port map( B1 => n1582_port, B2 => n11436, A => n11147, ZN 
                           => N2708);
   U16324 : OAI21_X1 port map( B1 => n1581_port, B2 => n11435, A => n11151, ZN 
                           => N2709);
   U16325 : OAI21_X1 port map( B1 => n1580_port, B2 => n11435, A => n11155, ZN 
                           => N2710);
   U16326 : OAI21_X1 port map( B1 => n1579_port, B2 => n11435, A => n11159, ZN 
                           => N2711);
   U16327 : OAI21_X1 port map( B1 => n1578_port, B2 => n11435, A => n11163, ZN 
                           => N2712);
   U16328 : OAI21_X1 port map( B1 => n1577_port, B2 => n11435, A => n11167, ZN 
                           => N2713);
   U16329 : OAI21_X1 port map( B1 => n1576_port, B2 => n11435, A => n11171, ZN 
                           => N2714);
   U16330 : OAI21_X1 port map( B1 => n1575_port, B2 => n11435, A => n11175, ZN 
                           => N2715);
   U16331 : OAI21_X1 port map( B1 => n1574_port, B2 => n11435, A => n11179, ZN 
                           => N2716);
   U16332 : OAI21_X1 port map( B1 => n1573_port, B2 => n11435, A => n11183, ZN 
                           => N2717);
   U16333 : OAI21_X1 port map( B1 => n1572_port, B2 => n11435, A => n11187, ZN 
                           => N2718);
   U16334 : OAI21_X1 port map( B1 => n1571_port, B2 => n11435, A => n11191, ZN 
                           => N2719);
   U16335 : OAI21_X1 port map( B1 => n1570_port, B2 => n11435, A => n11195, ZN 
                           => N2720);
   U16336 : OAI21_X1 port map( B1 => n1569_port, B2 => n11434, A => n11199, ZN 
                           => N2721);
   U16337 : OAI21_X1 port map( B1 => n1568_port, B2 => n11434, A => n11203, ZN 
                           => N2722);
   U16338 : OAI21_X1 port map( B1 => n1567_port, B2 => n11434, A => n11207, ZN 
                           => N2723);
   U16339 : OAI21_X1 port map( B1 => n1566_port, B2 => n11434, A => n11211, ZN 
                           => N2724);
   U16340 : OAI21_X1 port map( B1 => n1565_port, B2 => n11434, A => n11215, ZN 
                           => N2725);
   U16341 : OAI21_X1 port map( B1 => n1564_port, B2 => n11434, A => n11219, ZN 
                           => N2726);
   U16342 : OAI21_X1 port map( B1 => n1563_port, B2 => n11434, A => n11223, ZN 
                           => N2727);
   U16343 : OAI21_X1 port map( B1 => n1562_port, B2 => n11434, A => n11227, ZN 
                           => N2728);
   U16344 : OAI21_X1 port map( B1 => n1561_port, B2 => n11434, A => n11231, ZN 
                           => N2729);
   U16345 : OAI21_X1 port map( B1 => n1560_port, B2 => n11434, A => n11235, ZN 
                           => N2730);
   U16346 : OAI21_X1 port map( B1 => n1559_port, B2 => n11434, A => n11239, ZN 
                           => N2731);
   U16347 : OAI21_X1 port map( B1 => n1558_port, B2 => n11434, A => n11243, ZN 
                           => N2732);
   U16348 : OAI21_X1 port map( B1 => n1557_port, B2 => n11433, A => n11247, ZN 
                           => N2733);
   U16349 : OAI21_X1 port map( B1 => n1556_port, B2 => n11433, A => n11251, ZN 
                           => N2734);
   U16350 : OAI21_X1 port map( B1 => n1555_port, B2 => n11433, A => n11255, ZN 
                           => N2735);
   U16351 : OAI21_X1 port map( B1 => n1554_port, B2 => n11433, A => n11259, ZN 
                           => N2736);
   U16352 : OAI21_X1 port map( B1 => n1553_port, B2 => n11433, A => n11263, ZN 
                           => N2737);
   U16353 : OAI21_X1 port map( B1 => n1552_port, B2 => n11433, A => n11267, ZN 
                           => N2738);
   U16354 : OAI21_X1 port map( B1 => n1551_port, B2 => n11433, A => n11271, ZN 
                           => N2739);
   U16355 : OAI21_X1 port map( B1 => n1550_port, B2 => n11433, A => n11275, ZN 
                           => N2740);
   U16356 : OAI21_X1 port map( B1 => n1549_port, B2 => n11433, A => n11279, ZN 
                           => N2741);
   U16357 : OAI21_X1 port map( B1 => n1548_port, B2 => n11433, A => n11283, ZN 
                           => N2742);
   U16358 : OAI21_X1 port map( B1 => n1547_port, B2 => n11433, A => n11287, ZN 
                           => N2743);
   U16359 : OAI21_X1 port map( B1 => n1546_port, B2 => n11433, A => n11291, ZN 
                           => N2744);
   U16360 : OAI21_X1 port map( B1 => n1545_port, B2 => n11432, A => n11295, ZN 
                           => N2745);
   U16361 : OAI21_X1 port map( B1 => n1544_port, B2 => n11432, A => n11299, ZN 
                           => N2746);
   U16362 : OAI21_X1 port map( B1 => n1543_port, B2 => n11432, A => n11303, ZN 
                           => N2747);
   U16363 : OAI21_X1 port map( B1 => n1542_port, B2 => n11432, A => n11307, ZN 
                           => N2748);
   U16364 : OAI21_X1 port map( B1 => n1541_port, B2 => n11432, A => n11311, ZN 
                           => N2749);
   U16365 : OAI21_X1 port map( B1 => n1540_port, B2 => n11432, A => n11315, ZN 
                           => N2750);
   U16366 : OAI21_X1 port map( B1 => n1539_port, B2 => n11432, A => n11319, ZN 
                           => N2751);
   U16367 : OAI21_X1 port map( B1 => n1538_port, B2 => n11432, A => n11323, ZN 
                           => N2752);
   U16368 : OAI21_X1 port map( B1 => n1537_port, B2 => n11432, A => n11327, ZN 
                           => N2753);
   U16369 : OAI21_X1 port map( B1 => n1536_port, B2 => n11432, A => n11075, ZN 
                           => N2755);
   U16370 : OAI21_X1 port map( B1 => n1535_port, B2 => n11432, A => n11079, ZN 
                           => N2756);
   U16371 : OAI21_X1 port map( B1 => n1534_port, B2 => n11437, A => n11083, ZN 
                           => N2757);
   U16372 : OAI21_X1 port map( B1 => n1533_port, B2 => n11442, A => n11087, ZN 
                           => N2758);
   U16373 : OAI21_X1 port map( B1 => n1532_port, B2 => n11496, A => n11091, ZN 
                           => N2759);
   U16374 : OAI21_X1 port map( B1 => n1531_port, B2 => n11496, A => n11095, ZN 
                           => N2760);
   U16375 : OAI21_X1 port map( B1 => n1530_port, B2 => n11496, A => n11099, ZN 
                           => N2761);
   U16376 : OAI21_X1 port map( B1 => n1529_port, B2 => n11496, A => n11103, ZN 
                           => N2762);
   U16377 : OAI21_X1 port map( B1 => n1528_port, B2 => n11496, A => n11107, ZN 
                           => N2763);
   U16378 : OAI21_X1 port map( B1 => n1527_port, B2 => n11496, A => n11111, ZN 
                           => N2764);
   U16379 : OAI21_X1 port map( B1 => n1526_port, B2 => n11495, A => n11115, ZN 
                           => N2765);
   U16380 : OAI21_X1 port map( B1 => n1525_port, B2 => n11495, A => n11119, ZN 
                           => N2766);
   U16381 : OAI21_X1 port map( B1 => n1524_port, B2 => n11495, A => n11123, ZN 
                           => N2767);
   U16382 : OAI21_X1 port map( B1 => n1523_port, B2 => n11495, A => n11127, ZN 
                           => N2768);
   U16383 : OAI21_X1 port map( B1 => n1522_port, B2 => n11495, A => n11131, ZN 
                           => N2769);
   U16384 : OAI21_X1 port map( B1 => n1521_port, B2 => n11495, A => n11135, ZN 
                           => N2770);
   U16385 : OAI21_X1 port map( B1 => n1520_port, B2 => n11495, A => n11139, ZN 
                           => N2771);
   U16386 : OAI21_X1 port map( B1 => n1519_port, B2 => n11495, A => n11143, ZN 
                           => N2772);
   U16387 : OAI21_X1 port map( B1 => n1518_port, B2 => n11495, A => n11147, ZN 
                           => N2773);
   U16388 : OAI21_X1 port map( B1 => n1517_port, B2 => n11495, A => n11151, ZN 
                           => N2774);
   U16389 : OAI21_X1 port map( B1 => n1516_port, B2 => n11495, A => n11155, ZN 
                           => N2775);
   U16390 : OAI21_X1 port map( B1 => n1515_port, B2 => n11495, A => n11159, ZN 
                           => N2776);
   U16391 : OAI21_X1 port map( B1 => n1514_port, B2 => n11494, A => n11163, ZN 
                           => N2777);
   U16392 : OAI21_X1 port map( B1 => n1513_port, B2 => n11494, A => n11167, ZN 
                           => N2778);
   U16393 : OAI21_X1 port map( B1 => n1512_port, B2 => n11494, A => n11171, ZN 
                           => N2779);
   U16394 : OAI21_X1 port map( B1 => n1511_port, B2 => n11494, A => n11175, ZN 
                           => N2780);
   U16395 : OAI21_X1 port map( B1 => n1510_port, B2 => n11494, A => n11179, ZN 
                           => N2781);
   U16396 : OAI21_X1 port map( B1 => n1509_port, B2 => n11494, A => n11183, ZN 
                           => N2782);
   U16397 : OAI21_X1 port map( B1 => n1508_port, B2 => n11494, A => n11187, ZN 
                           => N2783);
   U16398 : OAI21_X1 port map( B1 => n1507_port, B2 => n11494, A => n11191, ZN 
                           => N2784);
   U16399 : OAI21_X1 port map( B1 => n1506_port, B2 => n11494, A => n11195, ZN 
                           => N2785);
   U16400 : OAI21_X1 port map( B1 => n1505_port, B2 => n11494, A => n11199, ZN 
                           => N2786);
   U16401 : OAI21_X1 port map( B1 => n1504_port, B2 => n11494, A => n11203, ZN 
                           => N2787);
   U16402 : OAI21_X1 port map( B1 => n1503_port, B2 => n11494, A => n11207, ZN 
                           => N2788);
   U16403 : OAI21_X1 port map( B1 => n1502_port, B2 => n11493, A => n11211, ZN 
                           => N2789);
   U16404 : OAI21_X1 port map( B1 => n1501_port, B2 => n11493, A => n11215, ZN 
                           => N2790);
   U16405 : OAI21_X1 port map( B1 => n1500_port, B2 => n11493, A => n11219, ZN 
                           => N2791);
   U16406 : OAI21_X1 port map( B1 => n1499_port, B2 => n11493, A => n11223, ZN 
                           => N2792);
   U16407 : OAI21_X1 port map( B1 => n1498_port, B2 => n11493, A => n11227, ZN 
                           => N2793);
   U16408 : OAI21_X1 port map( B1 => n1497_port, B2 => n11493, A => n11231, ZN 
                           => N2794);
   U16409 : OAI21_X1 port map( B1 => n1496_port, B2 => n11493, A => n11235, ZN 
                           => N2795);
   U16410 : OAI21_X1 port map( B1 => n1495_port, B2 => n11493, A => n11239, ZN 
                           => N2796);
   U16411 : OAI21_X1 port map( B1 => n1494_port, B2 => n11493, A => n11243, ZN 
                           => N2797);
   U16412 : OAI21_X1 port map( B1 => n1493_port, B2 => n11493, A => n11247, ZN 
                           => N2798);
   U16413 : OAI21_X1 port map( B1 => n1492_port, B2 => n11493, A => n11251, ZN 
                           => N2799);
   U16414 : OAI21_X1 port map( B1 => n1491_port, B2 => n11493, A => n11255, ZN 
                           => N2800);
   U16415 : OAI21_X1 port map( B1 => n1490_port, B2 => n11492, A => n11259, ZN 
                           => N2801);
   U16416 : OAI21_X1 port map( B1 => n1489_port, B2 => n11492, A => n11263, ZN 
                           => N2802);
   U16417 : OAI21_X1 port map( B1 => n1488_port, B2 => n11492, A => n11267, ZN 
                           => N2803);
   U16418 : OAI21_X1 port map( B1 => n1487_port, B2 => n11492, A => n11271, ZN 
                           => N2804);
   U16419 : OAI21_X1 port map( B1 => n1486_port, B2 => n11492, A => n11275, ZN 
                           => N2805);
   U16420 : OAI21_X1 port map( B1 => n1485_port, B2 => n11492, A => n11279, ZN 
                           => N2806);
   U16421 : OAI21_X1 port map( B1 => n1484_port, B2 => n11492, A => n11283, ZN 
                           => N2807);
   U16422 : OAI21_X1 port map( B1 => n1483_port, B2 => n11492, A => n11287, ZN 
                           => N2808);
   U16423 : OAI21_X1 port map( B1 => n1482_port, B2 => n11492, A => n11291, ZN 
                           => N2809);
   U16424 : OAI21_X1 port map( B1 => n1481_port, B2 => n11492, A => n11295, ZN 
                           => N2810);
   U16425 : OAI21_X1 port map( B1 => n1480_port, B2 => n11492, A => n11299, ZN 
                           => N2811);
   U16426 : OAI21_X1 port map( B1 => n1479_port, B2 => n11492, A => n11303, ZN 
                           => N2812);
   U16427 : OAI21_X1 port map( B1 => n1478_port, B2 => n11491, A => n11307, ZN 
                           => N2813);
   U16428 : OAI21_X1 port map( B1 => n1477_port, B2 => n11491, A => n11311, ZN 
                           => N2814);
   U16429 : OAI21_X1 port map( B1 => n1476_port, B2 => n11491, A => n11315, ZN 
                           => N2815);
   U16430 : OAI21_X1 port map( B1 => n1475_port, B2 => n11491, A => n11319, ZN 
                           => N2816);
   U16431 : OAI21_X1 port map( B1 => n1474_port, B2 => n11491, A => n11323, ZN 
                           => N2817);
   U16432 : OAI21_X1 port map( B1 => n1473_port, B2 => n11491, A => n11327, ZN 
                           => N2818);
   U16433 : OAI21_X1 port map( B1 => n1472_port, B2 => n11491, A => n11075, ZN 
                           => N2820);
   U16434 : OAI21_X1 port map( B1 => n1471_port, B2 => n11485, A => n11079, ZN 
                           => N2821);
   U16435 : OAI21_X1 port map( B1 => n1470_port, B2 => n11491, A => n11083, ZN 
                           => N2822);
   U16436 : OAI21_X1 port map( B1 => n1469_port, B2 => n11491, A => n11087, ZN 
                           => N2823);
   U16437 : OAI21_X1 port map( B1 => n1468_port, B2 => n11491, A => n11091, ZN 
                           => N2824);
   U16438 : OAI21_X1 port map( B1 => n1467_port, B2 => n11490, A => n11095, ZN 
                           => N2825);
   U16439 : OAI21_X1 port map( B1 => n1466_port, B2 => n11490, A => n11099, ZN 
                           => N2826);
   U16440 : OAI21_X1 port map( B1 => n1465_port, B2 => n11490, A => n11103, ZN 
                           => N2827);
   U16441 : OAI21_X1 port map( B1 => n1464_port, B2 => n11490, A => n11107, ZN 
                           => N2828);
   U16442 : OAI21_X1 port map( B1 => n1463_port, B2 => n11490, A => n11111, ZN 
                           => N2829);
   U16443 : OAI21_X1 port map( B1 => n1462_port, B2 => n11490, A => n11115, ZN 
                           => N2830);
   U16444 : OAI21_X1 port map( B1 => n1461_port, B2 => n11490, A => n11119, ZN 
                           => N2831);
   U16445 : OAI21_X1 port map( B1 => n1460_port, B2 => n11490, A => n11123, ZN 
                           => N2832);
   U16446 : OAI21_X1 port map( B1 => n1459_port, B2 => n11490, A => n11127, ZN 
                           => N2833);
   U16447 : OAI21_X1 port map( B1 => n1458_port, B2 => n11490, A => n11131, ZN 
                           => N2834);
   U16448 : OAI21_X1 port map( B1 => n1457_port, B2 => n11490, A => n11135, ZN 
                           => N2835);
   U16449 : OAI21_X1 port map( B1 => n1456_port, B2 => n11490, A => n11139, ZN 
                           => N2836);
   U16450 : OAI21_X1 port map( B1 => n1455_port, B2 => n11489, A => n11143, ZN 
                           => N2837);
   U16451 : OAI21_X1 port map( B1 => n1454_port, B2 => n11489, A => n11147, ZN 
                           => N2838);
   U16452 : OAI21_X1 port map( B1 => n1453_port, B2 => n11489, A => n11151, ZN 
                           => N2839);
   U16453 : OAI21_X1 port map( B1 => n1452_port, B2 => n11489, A => n11155, ZN 
                           => N2840);
   U16454 : OAI21_X1 port map( B1 => n1451_port, B2 => n11489, A => n11159, ZN 
                           => N2841);
   U16455 : OAI21_X1 port map( B1 => n1450_port, B2 => n11489, A => n11163, ZN 
                           => N2842);
   U16456 : OAI21_X1 port map( B1 => n1449_port, B2 => n11489, A => n11167, ZN 
                           => N2843);
   U16457 : OAI21_X1 port map( B1 => n1448_port, B2 => n11489, A => n11171, ZN 
                           => N2844);
   U16458 : OAI21_X1 port map( B1 => n1447_port, B2 => n11489, A => n11175, ZN 
                           => N2845);
   U16459 : OAI21_X1 port map( B1 => n1446_port, B2 => n11489, A => n11179, ZN 
                           => N2846);
   U16460 : OAI21_X1 port map( B1 => n1445_port, B2 => n11489, A => n11183, ZN 
                           => N2847);
   U16461 : OAI21_X1 port map( B1 => n1444_port, B2 => n11489, A => n11187, ZN 
                           => N2848);
   U16462 : OAI21_X1 port map( B1 => n1443_port, B2 => n11488, A => n11191, ZN 
                           => N2849);
   U16463 : OAI21_X1 port map( B1 => n1442_port, B2 => n11488, A => n11195, ZN 
                           => N2850);
   U16464 : OAI21_X1 port map( B1 => n1441_port, B2 => n11488, A => n11199, ZN 
                           => N2851);
   U16465 : OAI21_X1 port map( B1 => n1440_port, B2 => n11488, A => n11203, ZN 
                           => N2852);
   U16466 : OAI21_X1 port map( B1 => n1439_port, B2 => n11488, A => n11207, ZN 
                           => N2853);
   U16467 : OAI21_X1 port map( B1 => n1438_port, B2 => n11488, A => n11211, ZN 
                           => N2854);
   U16468 : OAI21_X1 port map( B1 => n1437_port, B2 => n11488, A => n11215, ZN 
                           => N2855);
   U16469 : OAI21_X1 port map( B1 => n1436_port, B2 => n11488, A => n11219, ZN 
                           => N2856);
   U16470 : OAI21_X1 port map( B1 => n1435_port, B2 => n11488, A => n11223, ZN 
                           => N2857);
   U16471 : OAI21_X1 port map( B1 => n1434_port, B2 => n11488, A => n11227, ZN 
                           => N2858);
   U16472 : OAI21_X1 port map( B1 => n1433_port, B2 => n11488, A => n11231, ZN 
                           => N2859);
   U16473 : OAI21_X1 port map( B1 => n1432_port, B2 => n11488, A => n11235, ZN 
                           => N2860);
   U16474 : OAI21_X1 port map( B1 => n1431_port, B2 => n11487, A => n11239, ZN 
                           => N2861);
   U16475 : OAI21_X1 port map( B1 => n1430_port, B2 => n11487, A => n11243, ZN 
                           => N2862);
   U16476 : OAI21_X1 port map( B1 => n1429_port, B2 => n11487, A => n11247, ZN 
                           => N2863);
   U16477 : OAI21_X1 port map( B1 => n1428_port, B2 => n11487, A => n11251, ZN 
                           => N2864);
   U16478 : OAI21_X1 port map( B1 => n1427_port, B2 => n11487, A => n11255, ZN 
                           => N2865);
   U16479 : OAI21_X1 port map( B1 => n1426_port, B2 => n11487, A => n11259, ZN 
                           => N2866);
   U16480 : OAI21_X1 port map( B1 => n1425_port, B2 => n11487, A => n11263, ZN 
                           => N2867);
   U16481 : OAI21_X1 port map( B1 => n1424_port, B2 => n11487, A => n11267, ZN 
                           => N2868);
   U16482 : OAI21_X1 port map( B1 => n1423_port, B2 => n11487, A => n11271, ZN 
                           => N2869);
   U16483 : OAI21_X1 port map( B1 => n1422_port, B2 => n11487, A => n11275, ZN 
                           => N2870);
   U16484 : OAI21_X1 port map( B1 => n1421_port, B2 => n11487, A => n11279, ZN 
                           => N2871);
   U16485 : OAI21_X1 port map( B1 => n1420_port, B2 => n11487, A => n11283, ZN 
                           => N2872);
   U16486 : OAI21_X1 port map( B1 => n1419_port, B2 => n11486, A => n11287, ZN 
                           => N2873);
   U16487 : OAI21_X1 port map( B1 => n1418_port, B2 => n11486, A => n11291, ZN 
                           => N2874);
   U16488 : OAI21_X1 port map( B1 => n1417_port, B2 => n11486, A => n11295, ZN 
                           => N2875);
   U16489 : OAI21_X1 port map( B1 => n1416_port, B2 => n11486, A => n11299, ZN 
                           => N2876);
   U16490 : OAI21_X1 port map( B1 => n1415_port, B2 => n11486, A => n11303, ZN 
                           => N2877);
   U16491 : OAI21_X1 port map( B1 => n1414_port, B2 => n11486, A => n11307, ZN 
                           => N2878);
   U16492 : OAI21_X1 port map( B1 => n1413_port, B2 => n11486, A => n11311, ZN 
                           => N2879);
   U16493 : OAI21_X1 port map( B1 => n1412_port, B2 => n11486, A => n11315, ZN 
                           => N2880);
   U16494 : OAI21_X1 port map( B1 => n1411_port, B2 => n11486, A => n11319, ZN 
                           => N2881);
   U16495 : OAI21_X1 port map( B1 => n1410_port, B2 => n11486, A => n11323, ZN 
                           => N2882);
   U16496 : OAI21_X1 port map( B1 => n1409_port, B2 => n11486, A => n11327, ZN 
                           => N2883);
   U16497 : OAI21_X1 port map( B1 => n1408_port, B2 => n11486, A => n11075, ZN 
                           => N2885);
   U16498 : OAI21_X1 port map( B1 => n1407_port, B2 => n11485, A => n11079, ZN 
                           => N2886);
   U16499 : OAI21_X1 port map( B1 => n1406_port, B2 => n11485, A => n11083, ZN 
                           => N2887);
   U16500 : OAI21_X1 port map( B1 => n1405_port, B2 => n11491, A => n11087, ZN 
                           => N2888);
   U16501 : OAI21_X1 port map( B1 => n1404_port, B2 => n11505, A => n11091, ZN 
                           => N2889);
   U16502 : OAI21_X1 port map( B1 => n1403_port, B2 => n11505, A => n11095, ZN 
                           => N2890);
   U16503 : OAI21_X1 port map( B1 => n1402_port, B2 => n11504, A => n11099, ZN 
                           => N2891);
   U16504 : OAI21_X1 port map( B1 => n1401_port, B2 => n11504, A => n11103, ZN 
                           => N2892);
   U16505 : OAI21_X1 port map( B1 => n1400_port, B2 => n11505, A => n11107, ZN 
                           => N2893);
   U16506 : OAI21_X1 port map( B1 => n1399_port, B2 => n11505, A => n11111, ZN 
                           => N2894);
   U16507 : OAI21_X1 port map( B1 => n1398_port, B2 => n11504, A => n11115, ZN 
                           => N2895);
   U16508 : OAI21_X1 port map( B1 => n1397_port, B2 => n11505, A => n11119, ZN 
                           => N2896);
   U16509 : OAI21_X1 port map( B1 => n1396_port, B2 => n11505, A => n11123, ZN 
                           => N2897);
   U16510 : OAI21_X1 port map( B1 => n1395_port, B2 => n11505, A => n11127, ZN 
                           => N2898);
   U16511 : OAI21_X1 port map( B1 => n1394_port, B2 => n11505, A => n11131, ZN 
                           => N2899);
   U16512 : OAI21_X1 port map( B1 => n1393_port, B2 => n11505, A => n11135, ZN 
                           => N2900);
   U16513 : OAI21_X1 port map( B1 => n1392_port, B2 => n11505, A => n11139, ZN 
                           => N2901);
   U16514 : OAI21_X1 port map( B1 => n1391_port, B2 => n11505, A => n11143, ZN 
                           => N2902);
   U16515 : OAI21_X1 port map( B1 => n1390_port, B2 => n11503, A => n11147, ZN 
                           => N2903);
   U16516 : OAI21_X1 port map( B1 => n1389_port, B2 => n11505, A => n11151, ZN 
                           => N2904);
   U16517 : OAI21_X1 port map( B1 => n1388_port, B2 => n11502, A => n11155, ZN 
                           => N2905);
   U16518 : OAI21_X1 port map( B1 => n1387_port, B2 => n11503, A => n11159, ZN 
                           => N2906);
   U16519 : OAI21_X1 port map( B1 => n1386_port, B2 => n11504, A => n11163, ZN 
                           => N2907);
   U16520 : OAI21_X1 port map( B1 => n1385_port, B2 => n11502, A => n11167, ZN 
                           => N2908);
   U16521 : OAI21_X1 port map( B1 => n1384_port, B2 => n11503, A => n11171, ZN 
                           => N2909);
   U16522 : OAI21_X1 port map( B1 => n1383_port, B2 => n11504, A => n11175, ZN 
                           => N2910);
   U16523 : OAI21_X1 port map( B1 => n1382_port, B2 => n11504, A => n11179, ZN 
                           => N2911);
   U16524 : OAI21_X1 port map( B1 => n1381_port, B2 => n11503, A => n11183, ZN 
                           => N2912);
   U16525 : OAI21_X1 port map( B1 => n1380_port, B2 => n11504, A => n11187, ZN 
                           => N2913);
   U16526 : OAI21_X1 port map( B1 => n1379_port, B2 => n11504, A => n11191, ZN 
                           => N2914);
   U16527 : OAI21_X1 port map( B1 => n1378_port, B2 => n11503, A => n11195, ZN 
                           => N2915);
   U16528 : OAI21_X1 port map( B1 => n1377_port, B2 => n11504, A => n11199, ZN 
                           => N2916);
   U16529 : OAI21_X1 port map( B1 => n1376_port, B2 => n11504, A => n11203, ZN 
                           => N2917);
   U16530 : OAI21_X1 port map( B1 => n1375_port, B2 => n11502, A => n11207, ZN 
                           => N2918);
   U16531 : OAI21_X1 port map( B1 => n1374_port, B2 => n11504, A => n11211, ZN 
                           => N2919);
   U16532 : OAI21_X1 port map( B1 => n1373_port, B2 => n11504, A => n11215, ZN 
                           => N2920);
   U16533 : OAI21_X1 port map( B1 => n1372_port, B2 => n11502, A => n11219, ZN 
                           => N2921);
   U16534 : OAI21_X1 port map( B1 => n1371_port, B2 => n11503, A => n11223, ZN 
                           => N2922);
   U16535 : OAI21_X1 port map( B1 => n1370_port, B2 => n11503, A => n11227, ZN 
                           => N2923);
   U16536 : OAI21_X1 port map( B1 => n1369_port, B2 => n11502, A => n11231, ZN 
                           => N2924);
   U16537 : OAI21_X1 port map( B1 => n1368_port, B2 => n11503, A => n11235, ZN 
                           => N2925);
   U16538 : OAI21_X1 port map( B1 => n1367_port, B2 => n11503, A => n11239, ZN 
                           => N2926);
   U16539 : OAI21_X1 port map( B1 => n1366_port, B2 => n11503, A => n11243, ZN 
                           => N2927);
   U16540 : OAI21_X1 port map( B1 => n1365_port, B2 => n11501, A => n11247, ZN 
                           => N2928);
   U16541 : OAI21_X1 port map( B1 => n1364_port, B2 => n11503, A => n11251, ZN 
                           => N2929);
   U16542 : OAI21_X1 port map( B1 => n1363_port, B2 => n11502, A => n11255, ZN 
                           => N2930);
   U16543 : OAI21_X1 port map( B1 => n1362_port, B2 => n11503, A => n11259, ZN 
                           => N2931);
   U16544 : OAI21_X1 port map( B1 => n1361_port, B2 => n11502, A => n11263, ZN 
                           => N2932);
   U16545 : OAI21_X1 port map( B1 => n1360_port, B2 => n11502, A => n11267, ZN 
                           => N2933);
   U16546 : OAI21_X1 port map( B1 => n1359_port, B2 => n11502, A => n11271, ZN 
                           => N2934);
   U16547 : OAI21_X1 port map( B1 => n1358_port, B2 => n11502, A => n11275, ZN 
                           => N2935);
   U16548 : OAI21_X1 port map( B1 => n1357_port, B2 => n11502, A => n11279, ZN 
                           => N2936);
   U16549 : OAI21_X1 port map( B1 => n1356_port, B2 => n11502, A => n11283, ZN 
                           => N2937);
   U16550 : OAI21_X1 port map( B1 => n1355_port, B2 => n11501, A => n11287, ZN 
                           => N2938);
   U16551 : OAI21_X1 port map( B1 => n1354_port, B2 => n11501, A => n11291, ZN 
                           => N2939);
   U16552 : OAI21_X1 port map( B1 => n1353_port, B2 => n11501, A => n11295, ZN 
                           => N2940);
   U16553 : OAI21_X1 port map( B1 => n1352_port, B2 => n11501, A => n11299, ZN 
                           => N2941);
   U16554 : OAI21_X1 port map( B1 => n1351_port, B2 => n11501, A => n11303, ZN 
                           => N2942);
   U16555 : OAI21_X1 port map( B1 => n1350_port, B2 => n11501, A => n11307, ZN 
                           => N2943);
   U16556 : OAI21_X1 port map( B1 => n1349_port, B2 => n11501, A => n11311, ZN 
                           => N2944);
   U16557 : OAI21_X1 port map( B1 => n1348_port, B2 => n11501, A => n11315, ZN 
                           => N2945);
   U16558 : OAI21_X1 port map( B1 => n1347_port, B2 => n11501, A => n11319, ZN 
                           => N2946);
   U16559 : OAI21_X1 port map( B1 => n1346_port, B2 => n11501, A => n11323, ZN 
                           => N2947);
   U16560 : OAI21_X1 port map( B1 => n1345_port, B2 => n11500, A => n11327, ZN 
                           => N2948);
   U16561 : OAI21_X1 port map( B1 => n1344_port, B2 => n11500, A => n11075, ZN 
                           => N2950);
   U16562 : OAI21_X1 port map( B1 => n1343_port, B2 => n11500, A => n11079, ZN 
                           => N2951);
   U16563 : OAI21_X1 port map( B1 => n1342_port, B2 => n11500, A => n11083, ZN 
                           => N2952);
   U16564 : OAI21_X1 port map( B1 => n1341_port, B2 => n11500, A => n11087, ZN 
                           => N2953);
   U16565 : OAI21_X1 port map( B1 => n1340_port, B2 => n11500, A => n11091, ZN 
                           => N2954);
   U16566 : OAI21_X1 port map( B1 => n1339_port, B2 => n11500, A => n11095, ZN 
                           => N2955);
   U16567 : OAI21_X1 port map( B1 => n1338_port, B2 => n11500, A => n11099, ZN 
                           => N2956);
   U16568 : OAI21_X1 port map( B1 => n1337_port, B2 => n11500, A => n11103, ZN 
                           => N2957);
   U16569 : OAI21_X1 port map( B1 => n1336_port, B2 => n11500, A => n11107, ZN 
                           => N2958);
   U16570 : OAI21_X1 port map( B1 => n1335_port, B2 => n11500, A => n11111, ZN 
                           => N2959);
   U16571 : OAI21_X1 port map( B1 => n1334_port, B2 => n11500, A => n11115, ZN 
                           => N2960);
   U16572 : OAI21_X1 port map( B1 => n1333_port, B2 => n11499, A => n11119, ZN 
                           => N2961);
   U16573 : OAI21_X1 port map( B1 => n1332_port, B2 => n11499, A => n11123, ZN 
                           => N2962);
   U16574 : OAI21_X1 port map( B1 => n1331_port, B2 => n11499, A => n11127, ZN 
                           => N2963);
   U16575 : OAI21_X1 port map( B1 => n1330_port, B2 => n11499, A => n11131, ZN 
                           => N2964);
   U16576 : OAI21_X1 port map( B1 => n1329_port, B2 => n11499, A => n11135, ZN 
                           => N2965);
   U16577 : OAI21_X1 port map( B1 => n1328_port, B2 => n11499, A => n11139, ZN 
                           => N2966);
   U16578 : OAI21_X1 port map( B1 => n1327_port, B2 => n11499, A => n11143, ZN 
                           => N2967);
   U16579 : OAI21_X1 port map( B1 => n1326_port, B2 => n11499, A => n11147, ZN 
                           => N2968);
   U16580 : OAI21_X1 port map( B1 => n1325_port, B2 => n11499, A => n11151, ZN 
                           => N2969);
   U16581 : OAI21_X1 port map( B1 => n1324_port, B2 => n11499, A => n11155, ZN 
                           => N2970);
   U16582 : OAI21_X1 port map( B1 => n1323_port, B2 => n11499, A => n11159, ZN 
                           => N2971);
   U16583 : OAI21_X1 port map( B1 => n1322_port, B2 => n11499, A => n11163, ZN 
                           => N2972);
   U16584 : OAI21_X1 port map( B1 => n1321_port, B2 => n11498, A => n11167, ZN 
                           => N2973);
   U16585 : OAI21_X1 port map( B1 => n1320_port, B2 => n11498, A => n11171, ZN 
                           => N2974);
   U16586 : OAI21_X1 port map( B1 => n1319_port, B2 => n11498, A => n11175, ZN 
                           => N2975);
   U16587 : OAI21_X1 port map( B1 => n1318_port, B2 => n11498, A => n11179, ZN 
                           => N2976);
   U16588 : OAI21_X1 port map( B1 => n1317_port, B2 => n11498, A => n11183, ZN 
                           => N2977);
   U16589 : OAI21_X1 port map( B1 => n1316_port, B2 => n11498, A => n11187, ZN 
                           => N2978);
   U16590 : OAI21_X1 port map( B1 => n1315_port, B2 => n11498, A => n11191, ZN 
                           => N2979);
   U16591 : OAI21_X1 port map( B1 => n1314_port, B2 => n11498, A => n11195, ZN 
                           => N2980);
   U16592 : OAI21_X1 port map( B1 => n1313_port, B2 => n11498, A => n11199, ZN 
                           => N2981);
   U16593 : OAI21_X1 port map( B1 => n1312_port, B2 => n11498, A => n11203, ZN 
                           => N2982);
   U16594 : OAI21_X1 port map( B1 => n1311_port, B2 => n11498, A => n11207, ZN 
                           => N2983);
   U16595 : OAI21_X1 port map( B1 => n1310_port, B2 => n11498, A => n11211, ZN 
                           => N2984);
   U16596 : OAI21_X1 port map( B1 => n1309_port, B2 => n11497, A => n11215, ZN 
                           => N2985);
   U16597 : OAI21_X1 port map( B1 => n1308_port, B2 => n11497, A => n11219, ZN 
                           => N2986);
   U16598 : OAI21_X1 port map( B1 => n1307_port, B2 => n11497, A => n11223, ZN 
                           => N2987);
   U16599 : OAI21_X1 port map( B1 => n1306_port, B2 => n11497, A => n11227, ZN 
                           => N2988);
   U16600 : OAI21_X1 port map( B1 => n1305_port, B2 => n11497, A => n11231, ZN 
                           => N2989);
   U16601 : OAI21_X1 port map( B1 => n1304_port, B2 => n11497, A => n11235, ZN 
                           => N2990);
   U16602 : OAI21_X1 port map( B1 => n1303_port, B2 => n11497, A => n11239, ZN 
                           => N2991);
   U16603 : OAI21_X1 port map( B1 => n1302_port, B2 => n11497, A => n11243, ZN 
                           => N2992);
   U16604 : OAI21_X1 port map( B1 => n1301_port, B2 => n11497, A => n11247, ZN 
                           => N2993);
   U16605 : OAI21_X1 port map( B1 => n1300_port, B2 => n11497, A => n11251, ZN 
                           => N2994);
   U16606 : OAI21_X1 port map( B1 => n1299_port, B2 => n11497, A => n11255, ZN 
                           => N2995);
   U16607 : OAI21_X1 port map( B1 => n1298_port, B2 => n11497, A => n11259, ZN 
                           => N2996);
   U16608 : OAI21_X1 port map( B1 => n1297_port, B2 => n11496, A => n11263, ZN 
                           => N2997);
   U16609 : OAI21_X1 port map( B1 => n1296_port, B2 => n11496, A => n11267, ZN 
                           => N2998);
   U16610 : OAI21_X1 port map( B1 => n1295_port, B2 => n11496, A => n11271, ZN 
                           => N2999);
   U16611 : OAI21_X1 port map( B1 => n1294_port, B2 => n11496, A => n11275, ZN 
                           => N3000);
   U16612 : OAI21_X1 port map( B1 => n1293_port, B2 => n11496, A => n11279, ZN 
                           => N3001);
   U16613 : OAI21_X1 port map( B1 => n1292_port, B2 => n11496, A => n11283, ZN 
                           => N3002);
   U16614 : OAI21_X1 port map( B1 => n1291_port, B2 => n11501, A => n11287, ZN 
                           => N3003);
   U16615 : OAI21_X1 port map( B1 => n1290_port, B2 => n11475, A => n11291, ZN 
                           => N3004);
   U16616 : OAI21_X1 port map( B1 => n1289_port, B2 => n11474, A => n11295, ZN 
                           => N3005);
   U16617 : OAI21_X1 port map( B1 => n1288_port, B2 => n11474, A => n11299, ZN 
                           => N3006);
   U16618 : OAI21_X1 port map( B1 => n1287_port, B2 => n11474, A => n11303, ZN 
                           => N3007);
   U16619 : OAI21_X1 port map( B1 => n1286_port, B2 => n11474, A => n11307, ZN 
                           => N3008);
   U16620 : OAI21_X1 port map( B1 => n1285_port, B2 => n11474, A => n11311, ZN 
                           => N3009);
   U16621 : OAI21_X1 port map( B1 => n1284_port, B2 => n11474, A => n11315, ZN 
                           => N3010);
   U16622 : OAI21_X1 port map( B1 => n1283_port, B2 => n11474, A => n11319, ZN 
                           => N3011);
   U16623 : OAI21_X1 port map( B1 => n1282_port, B2 => n11474, A => n11323, ZN 
                           => N3012);
   U16624 : OAI21_X1 port map( B1 => n1281_port, B2 => n11474, A => n11327, ZN 
                           => N3013);
   U16625 : OAI21_X1 port map( B1 => n1280_port, B2 => n11474, A => n11076, ZN 
                           => N3015);
   U16626 : OAI21_X1 port map( B1 => n1279_port, B2 => n11474, A => n11080, ZN 
                           => N3016);
   U16627 : OAI21_X1 port map( B1 => n1278_port, B2 => n11474, A => n11084, ZN 
                           => N3017);
   U16628 : OAI21_X1 port map( B1 => n1277_port, B2 => n11473, A => n11088, ZN 
                           => N3018);
   U16629 : OAI21_X1 port map( B1 => n1276_port, B2 => n11473, A => n11092, ZN 
                           => N3019);
   U16630 : OAI21_X1 port map( B1 => n1275_port, B2 => n11473, A => n11096, ZN 
                           => N3020);
   U16631 : OAI21_X1 port map( B1 => n1274_port, B2 => n11473, A => n11100, ZN 
                           => N3021);
   U16632 : OAI21_X1 port map( B1 => n1273_port, B2 => n11473, A => n11104, ZN 
                           => N3022);
   U16633 : OAI21_X1 port map( B1 => n1272_port, B2 => n11473, A => n11108, ZN 
                           => N3023);
   U16634 : OAI21_X1 port map( B1 => n1271_port, B2 => n11473, A => n11112, ZN 
                           => N3024);
   U16635 : OAI21_X1 port map( B1 => n1270_port, B2 => n11473, A => n11116, ZN 
                           => N3025);
   U16636 : OAI21_X1 port map( B1 => n1269_port, B2 => n11473, A => n11120, ZN 
                           => N3026);
   U16637 : OAI21_X1 port map( B1 => n1268_port, B2 => n11473, A => n11124, ZN 
                           => N3027);
   U16638 : OAI21_X1 port map( B1 => n1267_port, B2 => n11473, A => n11128, ZN 
                           => N3028);
   U16639 : OAI21_X1 port map( B1 => n1266_port, B2 => n11473, A => n11132, ZN 
                           => N3029);
   U16640 : OAI21_X1 port map( B1 => n1265_port, B2 => n11472, A => n11136, ZN 
                           => N3030);
   U16641 : OAI21_X1 port map( B1 => n1264_port, B2 => n11472, A => n11140, ZN 
                           => N3031);
   U16642 : OAI21_X1 port map( B1 => n1263_port, B2 => n11472, A => n11144, ZN 
                           => N3032);
   U16643 : OAI21_X1 port map( B1 => n1262_port, B2 => n11472, A => n11148, ZN 
                           => N3033);
   U16644 : OAI21_X1 port map( B1 => n1261_port, B2 => n11472, A => n11152, ZN 
                           => N3034);
   U16645 : OAI21_X1 port map( B1 => n1260_port, B2 => n11472, A => n11156, ZN 
                           => N3035);
   U16646 : OAI21_X1 port map( B1 => n1259_port, B2 => n11472, A => n11160, ZN 
                           => N3036);
   U16647 : OAI21_X1 port map( B1 => n1258_port, B2 => n11472, A => n11164, ZN 
                           => N3037);
   U16648 : OAI21_X1 port map( B1 => n1257_port, B2 => n11472, A => n11168, ZN 
                           => N3038);
   U16649 : OAI21_X1 port map( B1 => n1256_port, B2 => n11472, A => n11172, ZN 
                           => N3039);
   U16650 : OAI21_X1 port map( B1 => n1255_port, B2 => n11472, A => n11176, ZN 
                           => N3040);
   U16651 : OAI21_X1 port map( B1 => n1254_port, B2 => n11472, A => n11180, ZN 
                           => N3041);
   U16652 : OAI21_X1 port map( B1 => n1253_port, B2 => n11471, A => n11184, ZN 
                           => N3042);
   U16653 : OAI21_X1 port map( B1 => n1252_port, B2 => n11471, A => n11188, ZN 
                           => N3043);
   U16654 : OAI21_X1 port map( B1 => n1251_port, B2 => n11471, A => n11192, ZN 
                           => N3044);
   U16655 : OAI21_X1 port map( B1 => n1250_port, B2 => n11471, A => n11196, ZN 
                           => N3045);
   U16656 : OAI21_X1 port map( B1 => n1249_port, B2 => n11471, A => n11200, ZN 
                           => N3046);
   U16657 : OAI21_X1 port map( B1 => n1248_port, B2 => n11471, A => n11204, ZN 
                           => N3047);
   U16658 : OAI21_X1 port map( B1 => n1247_port, B2 => n11471, A => n11208, ZN 
                           => N3048);
   U16659 : OAI21_X1 port map( B1 => n1246_port, B2 => n11471, A => n11212, ZN 
                           => N3049);
   U16660 : OAI21_X1 port map( B1 => n1245_port, B2 => n11471, A => n11216, ZN 
                           => N3050);
   U16661 : OAI21_X1 port map( B1 => n1244_port, B2 => n11471, A => n11220, ZN 
                           => N3051);
   U16662 : OAI21_X1 port map( B1 => n1243_port, B2 => n11471, A => n11224, ZN 
                           => N3052);
   U16663 : OAI21_X1 port map( B1 => n1242_port, B2 => n11471, A => n11228, ZN 
                           => N3053);
   U16664 : OAI21_X1 port map( B1 => n1241_port, B2 => n11470, A => n11232, ZN 
                           => N3054);
   U16665 : OAI21_X1 port map( B1 => n1240_port, B2 => n11470, A => n11236, ZN 
                           => N3055);
   U16666 : OAI21_X1 port map( B1 => n1239_port, B2 => n11470, A => n11240, ZN 
                           => N3056);
   U16667 : OAI21_X1 port map( B1 => n1238_port, B2 => n11470, A => n11244, ZN 
                           => N3057);
   U16668 : OAI21_X1 port map( B1 => n1237_port, B2 => n11470, A => n11248, ZN 
                           => N3058);
   U16669 : OAI21_X1 port map( B1 => n1236_port, B2 => n11470, A => n11252, ZN 
                           => N3059);
   U16670 : OAI21_X1 port map( B1 => n1235_port, B2 => n11470, A => n11256, ZN 
                           => N3060);
   U16671 : OAI21_X1 port map( B1 => n1234_port, B2 => n11470, A => n11260, ZN 
                           => N3061);
   U16672 : OAI21_X1 port map( B1 => n1233_port, B2 => n11470, A => n11264, ZN 
                           => N3062);
   U16673 : OAI21_X1 port map( B1 => n1232_port, B2 => n11470, A => n11268, ZN 
                           => N3063);
   U16674 : OAI21_X1 port map( B1 => n1231_port, B2 => n11470, A => n11272, ZN 
                           => N3064);
   U16675 : OAI21_X1 port map( B1 => n1230_port, B2 => n11470, A => n11276, ZN 
                           => N3065);
   U16676 : OAI21_X1 port map( B1 => n1229_port, B2 => n11469, A => n11280, ZN 
                           => N3066);
   U16677 : OAI21_X1 port map( B1 => n1228_port, B2 => n11469, A => n11284, ZN 
                           => N3067);
   U16678 : OAI21_X1 port map( B1 => n1227_port, B2 => n11469, A => n11288, ZN 
                           => N3068);
   U16679 : OAI21_X1 port map( B1 => n1226_port, B2 => n11469, A => n11292, ZN 
                           => N3069);
   U16680 : OAI21_X1 port map( B1 => n1225_port, B2 => n11469, A => n11296, ZN 
                           => N3070);
   U16681 : OAI21_X1 port map( B1 => n1224_port, B2 => n11469, A => n11300, ZN 
                           => N3071);
   U16682 : OAI21_X1 port map( B1 => n1223_port, B2 => n11469, A => n11304, ZN 
                           => N3072);
   U16683 : OAI21_X1 port map( B1 => n1222_port, B2 => n11469, A => n11308, ZN 
                           => N3073);
   U16684 : OAI21_X1 port map( B1 => n1221_port, B2 => n11469, A => n11312, ZN 
                           => N3074);
   U16685 : OAI21_X1 port map( B1 => n1220_port, B2 => n11469, A => n11316, ZN 
                           => N3075);
   U16686 : OAI21_X1 port map( B1 => n1219_port, B2 => n11469, A => n11320, ZN 
                           => N3076);
   U16687 : OAI21_X1 port map( B1 => n1218_port, B2 => n11468, A => n11324, ZN 
                           => N3077);
   U16688 : OAI21_X1 port map( B1 => n1217_port, B2 => n11468, A => n11328, ZN 
                           => N3078);
   U16689 : OAI21_X1 port map( B1 => n1216_port, B2 => n11468, A => n11076, ZN 
                           => N3080);
   U16690 : OAI21_X1 port map( B1 => n1215_port, B2 => n11468, A => n11080, ZN 
                           => N3081);
   U16691 : OAI21_X1 port map( B1 => n1214_port, B2 => n11468, A => n11084, ZN 
                           => N3082);
   U16692 : OAI21_X1 port map( B1 => n1213_port, B2 => n11468, A => n11088, ZN 
                           => N3083);
   U16693 : OAI21_X1 port map( B1 => n1212_port, B2 => n11468, A => n11092, ZN 
                           => N3084);
   U16694 : OAI21_X1 port map( B1 => n1211_port, B2 => n11468, A => n11096, ZN 
                           => N3085);
   U16695 : OAI21_X1 port map( B1 => n1210_port, B2 => n11468, A => n11100, ZN 
                           => N3086);
   U16696 : OAI21_X1 port map( B1 => n1209_port, B2 => n11468, A => n11104, ZN 
                           => N3087);
   U16697 : OAI21_X1 port map( B1 => n1208_port, B2 => n11468, A => n11108, ZN 
                           => N3088);
   U16698 : OAI21_X1 port map( B1 => n1207_port, B2 => n11468, A => n11112, ZN 
                           => N3089);
   U16699 : OAI21_X1 port map( B1 => n1206_port, B2 => n11467, A => n11116, ZN 
                           => N3090);
   U16700 : OAI21_X1 port map( B1 => n1205_port, B2 => n11467, A => n11120, ZN 
                           => N3091);
   U16701 : OAI21_X1 port map( B1 => n1204_port, B2 => n11467, A => n11124, ZN 
                           => N3092);
   U16702 : OAI21_X1 port map( B1 => n1203_port, B2 => n11467, A => n11128, ZN 
                           => N3093);
   U16703 : OAI21_X1 port map( B1 => n1202_port, B2 => n11467, A => n11132, ZN 
                           => N3094);
   U16704 : OAI21_X1 port map( B1 => n1201_port, B2 => n11467, A => n11136, ZN 
                           => N3095);
   U16705 : OAI21_X1 port map( B1 => n1200_port, B2 => n11467, A => n11140, ZN 
                           => N3096);
   U16706 : OAI21_X1 port map( B1 => n1199_port, B2 => n11467, A => n11144, ZN 
                           => N3097);
   U16707 : OAI21_X1 port map( B1 => n1198_port, B2 => n11467, A => n11148, ZN 
                           => N3098);
   U16708 : OAI21_X1 port map( B1 => n1197_port, B2 => n11467, A => n11152, ZN 
                           => N3099);
   U16709 : OAI21_X1 port map( B1 => n1196_port, B2 => n11467, A => n11156, ZN 
                           => N3100);
   U16710 : OAI21_X1 port map( B1 => n1195_port, B2 => n11467, A => n11160, ZN 
                           => N3101);
   U16711 : OAI21_X1 port map( B1 => n1194_port, B2 => n11466, A => n11164, ZN 
                           => N3102);
   U16712 : OAI21_X1 port map( B1 => n1193_port, B2 => n11466, A => n11168, ZN 
                           => N3103);
   U16713 : OAI21_X1 port map( B1 => n1192_port, B2 => n11466, A => n11172, ZN 
                           => N3104);
   U16714 : OAI21_X1 port map( B1 => n1191_port, B2 => n11466, A => n11176, ZN 
                           => N3105);
   U16715 : OAI21_X1 port map( B1 => n1190_port, B2 => n11466, A => n11180, ZN 
                           => N3106);
   U16716 : OAI21_X1 port map( B1 => n1189_port, B2 => n11466, A => n11184, ZN 
                           => N3107);
   U16717 : OAI21_X1 port map( B1 => n1188_port, B2 => n11466, A => n11188, ZN 
                           => N3108);
   U16718 : OAI21_X1 port map( B1 => n1187_port, B2 => n11466, A => n11192, ZN 
                           => N3109);
   U16719 : OAI21_X1 port map( B1 => n1186_port, B2 => n11466, A => n11196, ZN 
                           => N3110);
   U16720 : OAI21_X1 port map( B1 => n1185_port, B2 => n11466, A => n11200, ZN 
                           => N3111);
   U16721 : OAI21_X1 port map( B1 => n1184_port, B2 => n11466, A => n11204, ZN 
                           => N3112);
   U16722 : OAI21_X1 port map( B1 => n1183_port, B2 => n11466, A => n11208, ZN 
                           => N3113);
   U16723 : OAI21_X1 port map( B1 => n1182_port, B2 => n11465, A => n11212, ZN 
                           => N3114);
   U16724 : OAI21_X1 port map( B1 => n1181_port, B2 => n11465, A => n11216, ZN 
                           => N3115);
   U16725 : OAI21_X1 port map( B1 => n1180_port, B2 => n11465, A => n11220, ZN 
                           => N3116);
   U16726 : OAI21_X1 port map( B1 => n1179_port, B2 => n11465, A => n11224, ZN 
                           => N3117);
   U16727 : OAI21_X1 port map( B1 => n1178_port, B2 => n11465, A => n11228, ZN 
                           => N3118);
   U16728 : OAI21_X1 port map( B1 => n1177_port, B2 => n11465, A => n11232, ZN 
                           => N3119);
   U16729 : OAI21_X1 port map( B1 => n1176_port, B2 => n11465, A => n11236, ZN 
                           => N3120);
   U16730 : OAI21_X1 port map( B1 => n1175_port, B2 => n11465, A => n11240, ZN 
                           => N3121);
   U16731 : OAI21_X1 port map( B1 => n1174_port, B2 => n11465, A => n11244, ZN 
                           => N3122);
   U16732 : OAI21_X1 port map( B1 => n1173_port, B2 => n11465, A => n11248, ZN 
                           => N3123);
   U16733 : OAI21_X1 port map( B1 => n1172_port, B2 => n11465, A => n11252, ZN 
                           => N3124);
   U16734 : OAI21_X1 port map( B1 => n1171_port, B2 => n11465, A => n11256, ZN 
                           => N3125);
   U16735 : OAI21_X1 port map( B1 => n1170_port, B2 => n11464, A => n11260, ZN 
                           => N3126);
   U16736 : OAI21_X1 port map( B1 => n1169_port, B2 => n11464, A => n11264, ZN 
                           => N3127);
   U16737 : OAI21_X1 port map( B1 => n1168_port, B2 => n11464, A => n11268, ZN 
                           => N3128);
   U16738 : OAI21_X1 port map( B1 => n1167_port, B2 => n11464, A => n11272, ZN 
                           => N3129);
   U16739 : OAI21_X1 port map( B1 => n1166_port, B2 => n11464, A => n11276, ZN 
                           => N3130);
   U16740 : OAI21_X1 port map( B1 => n1165_port, B2 => n11464, A => n11280, ZN 
                           => N3131);
   U16741 : OAI21_X1 port map( B1 => n1164_port, B2 => n11464, A => n11284, ZN 
                           => N3132);
   U16742 : OAI21_X1 port map( B1 => n1163_port, B2 => n11464, A => n11288, ZN 
                           => N3133);
   U16743 : OAI21_X1 port map( B1 => n1162_port, B2 => n11469, A => n11292, ZN 
                           => N3134);
   U16744 : OAI21_X1 port map( B1 => n1161_port, B2 => n11485, A => n11296, ZN 
                           => N3135);
   U16745 : OAI21_X1 port map( B1 => n1160_port, B2 => n11485, A => n11300, ZN 
                           => N3136);
   U16746 : OAI21_X1 port map( B1 => n1159_port, B2 => n11485, A => n11304, ZN 
                           => N3137);
   U16747 : OAI21_X1 port map( B1 => n1158_port, B2 => n11485, A => n11308, ZN 
                           => N3138);
   U16748 : OAI21_X1 port map( B1 => n1157_port, B2 => n11485, A => n11312, ZN 
                           => N3139);
   U16749 : OAI21_X1 port map( B1 => n1156_port, B2 => n11485, A => n11316, ZN 
                           => N3140);
   U16750 : OAI21_X1 port map( B1 => n1155_port, B2 => n11485, A => n11320, ZN 
                           => N3141);
   U16751 : OAI21_X1 port map( B1 => n1154_port, B2 => n11485, A => n11324, ZN 
                           => N3142);
   U16752 : OAI21_X1 port map( B1 => n1153_port, B2 => n11485, A => n11328, ZN 
                           => N3143);
   U16753 : OAI21_X1 port map( B1 => n1152_port, B2 => n11484, A => n11076, ZN 
                           => N3145);
   U16754 : OAI21_X1 port map( B1 => n1151_port, B2 => n11484, A => n11080, ZN 
                           => N3146);
   U16755 : OAI21_X1 port map( B1 => n1150_port, B2 => n11484, A => n11084, ZN 
                           => N3147);
   U16756 : OAI21_X1 port map( B1 => n1149_port, B2 => n11484, A => n11088, ZN 
                           => N3148);
   U16757 : OAI21_X1 port map( B1 => n1148_port, B2 => n11484, A => n11092, ZN 
                           => N3149);
   U16758 : OAI21_X1 port map( B1 => n1147_port, B2 => n11484, A => n11096, ZN 
                           => N3150);
   U16759 : OAI21_X1 port map( B1 => n1146_port, B2 => n11484, A => n11100, ZN 
                           => N3151);
   U16760 : OAI21_X1 port map( B1 => n1145_port, B2 => n11484, A => n11104, ZN 
                           => N3152);
   U16761 : OAI21_X1 port map( B1 => n1144_port, B2 => n11484, A => n11108, ZN 
                           => N3153);
   U16762 : OAI21_X1 port map( B1 => n1143_port, B2 => n11484, A => n11112, ZN 
                           => N3154);
   U16763 : OAI21_X1 port map( B1 => n1142_port, B2 => n11484, A => n11116, ZN 
                           => N3155);
   U16764 : OAI21_X1 port map( B1 => n1141_port, B2 => n11484, A => n11120, ZN 
                           => N3156);
   U16765 : OAI21_X1 port map( B1 => n1140_port, B2 => n11483, A => n11124, ZN 
                           => N3157);
   U16766 : OAI21_X1 port map( B1 => n1139_port, B2 => n11483, A => n11128, ZN 
                           => N3158);
   U16767 : OAI21_X1 port map( B1 => n1138_port, B2 => n11483, A => n11132, ZN 
                           => N3159);
   U16768 : OAI21_X1 port map( B1 => n1137_port, B2 => n11483, A => n11136, ZN 
                           => N3160);
   U16769 : OAI21_X1 port map( B1 => n1136_port, B2 => n11483, A => n11140, ZN 
                           => N3161);
   U16770 : OAI21_X1 port map( B1 => n1135_port, B2 => n11483, A => n11144, ZN 
                           => N3162);
   U16771 : OAI21_X1 port map( B1 => n1134_port, B2 => n11483, A => n11148, ZN 
                           => N3163);
   U16772 : OAI21_X1 port map( B1 => n1133_port, B2 => n11483, A => n11152, ZN 
                           => N3164);
   U16773 : OAI21_X1 port map( B1 => n1132_port, B2 => n11483, A => n11156, ZN 
                           => N3165);
   U16774 : OAI21_X1 port map( B1 => n1131_port, B2 => n11483, A => n11160, ZN 
                           => N3166);
   U16775 : OAI21_X1 port map( B1 => n1130_port, B2 => n11483, A => n11164, ZN 
                           => N3167);
   U16776 : OAI21_X1 port map( B1 => n1129_port, B2 => n11483, A => n11168, ZN 
                           => N3168);
   U16777 : OAI21_X1 port map( B1 => n1128_port, B2 => n11482, A => n11172, ZN 
                           => N3169);
   U16778 : OAI21_X1 port map( B1 => n1127_port, B2 => n11482, A => n11176, ZN 
                           => N3170);
   U16779 : OAI21_X1 port map( B1 => n1126_port, B2 => n11482, A => n11180, ZN 
                           => N3171);
   U16780 : OAI21_X1 port map( B1 => n1125_port, B2 => n11482, A => n11184, ZN 
                           => N3172);
   U16781 : OAI21_X1 port map( B1 => n1124_port, B2 => n11482, A => n11188, ZN 
                           => N3173);
   U16782 : OAI21_X1 port map( B1 => n1123_port, B2 => n11482, A => n11192, ZN 
                           => N3174);
   U16783 : OAI21_X1 port map( B1 => n1122_port, B2 => n11482, A => n11196, ZN 
                           => N3175);
   U16784 : OAI21_X1 port map( B1 => n1121_port, B2 => n11482, A => n11200, ZN 
                           => N3176);
   U16785 : OAI21_X1 port map( B1 => n1120_port, B2 => n11482, A => n11204, ZN 
                           => N3177);
   U16786 : OAI21_X1 port map( B1 => n1119_port, B2 => n11482, A => n11208, ZN 
                           => N3178);
   U16787 : OAI21_X1 port map( B1 => n1118_port, B2 => n11482, A => n11212, ZN 
                           => N3179);
   U16788 : OAI21_X1 port map( B1 => n1117_port, B2 => n11482, A => n11216, ZN 
                           => N3180);
   U16789 : OAI21_X1 port map( B1 => n1116_port, B2 => n11481, A => n11220, ZN 
                           => N3181);
   U16790 : OAI21_X1 port map( B1 => n1115_port, B2 => n11481, A => n11224, ZN 
                           => N3182);
   U16791 : OAI21_X1 port map( B1 => n1114_port, B2 => n11481, A => n11228, ZN 
                           => N3183);
   U16792 : OAI21_X1 port map( B1 => n1113_port, B2 => n11481, A => n11232, ZN 
                           => N3184);
   U16793 : OAI21_X1 port map( B1 => n1112_port, B2 => n11481, A => n11236, ZN 
                           => N3185);
   U16794 : OAI21_X1 port map( B1 => n1111_port, B2 => n11481, A => n11240, ZN 
                           => N3186);
   U16795 : OAI21_X1 port map( B1 => n1110_port, B2 => n11481, A => n11244, ZN 
                           => N3187);
   U16796 : OAI21_X1 port map( B1 => n1109_port, B2 => n11481, A => n11248, ZN 
                           => N3188);
   U16797 : OAI21_X1 port map( B1 => n1108_port, B2 => n11481, A => n11252, ZN 
                           => N3189);
   U16798 : OAI21_X1 port map( B1 => n1107_port, B2 => n11481, A => n11256, ZN 
                           => N3190);
   U16799 : OAI21_X1 port map( B1 => n1106_port, B2 => n11481, A => n11260, ZN 
                           => N3191);
   U16800 : OAI21_X1 port map( B1 => n1105_port, B2 => n11481, A => n11264, ZN 
                           => N3192);
   U16801 : OAI21_X1 port map( B1 => n1104_port, B2 => n11480, A => n11268, ZN 
                           => N3193);
   U16802 : OAI21_X1 port map( B1 => n1103_port, B2 => n11480, A => n11272, ZN 
                           => N3194);
   U16803 : OAI21_X1 port map( B1 => n1102_port, B2 => n11480, A => n11276, ZN 
                           => N3195);
   U16804 : OAI21_X1 port map( B1 => n1101_port, B2 => n11480, A => n11280, ZN 
                           => N3196);
   U16805 : OAI21_X1 port map( B1 => n1100_port, B2 => n11480, A => n11284, ZN 
                           => N3197);
   U16806 : OAI21_X1 port map( B1 => n1099_port, B2 => n11480, A => n11288, ZN 
                           => N3198);
   U16807 : OAI21_X1 port map( B1 => n1098_port, B2 => n11480, A => n11292, ZN 
                           => N3199);
   U16808 : OAI21_X1 port map( B1 => n1097_port, B2 => n11480, A => n11296, ZN 
                           => N3200);
   U16809 : OAI21_X1 port map( B1 => n1096_port, B2 => n11480, A => n11300, ZN 
                           => N3201);
   U16810 : OAI21_X1 port map( B1 => n1095_port, B2 => n11480, A => n11304, ZN 
                           => N3202);
   U16811 : OAI21_X1 port map( B1 => n1094_port, B2 => n11480, A => n11308, ZN 
                           => N3203);
   U16812 : OAI21_X1 port map( B1 => n1093_port, B2 => n11479, A => n11312, ZN 
                           => N3204);
   U16813 : OAI21_X1 port map( B1 => n1092_port, B2 => n11479, A => n11316, ZN 
                           => N3205);
   U16814 : OAI21_X1 port map( B1 => n1091_port, B2 => n11479, A => n11320, ZN 
                           => N3206);
   U16815 : OAI21_X1 port map( B1 => n1090_port, B2 => n11479, A => n11324, ZN 
                           => N3207);
   U16816 : OAI21_X1 port map( B1 => n1089_port, B2 => n11479, A => n11328, ZN 
                           => N3208);
   U16817 : OAI21_X1 port map( B1 => n1088_port, B2 => n11479, A => n11076, ZN 
                           => N3210);
   U16818 : OAI21_X1 port map( B1 => n1087_port, B2 => n11479, A => n11080, ZN 
                           => N3211);
   U16819 : OAI21_X1 port map( B1 => n1086_port, B2 => n11479, A => n11084, ZN 
                           => N3212);
   U16820 : OAI21_X1 port map( B1 => n1085_port, B2 => n11479, A => n11088, ZN 
                           => N3213);
   U16821 : OAI21_X1 port map( B1 => n1084_port, B2 => n11479, A => n11092, ZN 
                           => N3214);
   U16822 : OAI21_X1 port map( B1 => n1083_port, B2 => n11479, A => n11096, ZN 
                           => N3215);
   U16823 : OAI21_X1 port map( B1 => n1082_port, B2 => n11479, A => n11100, ZN 
                           => N3216);
   U16824 : OAI21_X1 port map( B1 => n1081_port, B2 => n11478, A => n11104, ZN 
                           => N3217);
   U16825 : OAI21_X1 port map( B1 => n1080_port, B2 => n11478, A => n11108, ZN 
                           => N3218);
   U16826 : OAI21_X1 port map( B1 => n1079_port, B2 => n11478, A => n11112, ZN 
                           => N3219);
   U16827 : OAI21_X1 port map( B1 => n1078_port, B2 => n11478, A => n11116, ZN 
                           => N3220);
   U16828 : OAI21_X1 port map( B1 => n1077_port, B2 => n11478, A => n11120, ZN 
                           => N3221);
   U16829 : OAI21_X1 port map( B1 => n1076_port, B2 => n11478, A => n11124, ZN 
                           => N3222);
   U16830 : OAI21_X1 port map( B1 => n1075_port, B2 => n11478, A => n11128, ZN 
                           => N3223);
   U16831 : OAI21_X1 port map( B1 => n1074_port, B2 => n11478, A => n11132, ZN 
                           => N3224);
   U16832 : OAI21_X1 port map( B1 => n1073_port, B2 => n11478, A => n11136, ZN 
                           => N3225);
   U16833 : OAI21_X1 port map( B1 => n1072_port, B2 => n11478, A => n11140, ZN 
                           => N3226);
   U16834 : OAI21_X1 port map( B1 => n1071_port, B2 => n11478, A => n11144, ZN 
                           => N3227);
   U16835 : OAI21_X1 port map( B1 => n1070_port, B2 => n11478, A => n11148, ZN 
                           => N3228);
   U16836 : OAI21_X1 port map( B1 => n1069_port, B2 => n11477, A => n11152, ZN 
                           => N3229);
   U16837 : OAI21_X1 port map( B1 => n1068_port, B2 => n11477, A => n11156, ZN 
                           => N3230);
   U16838 : OAI21_X1 port map( B1 => n1067_port, B2 => n11477, A => n11160, ZN 
                           => N3231);
   U16839 : OAI21_X1 port map( B1 => n1066_port, B2 => n11477, A => n11164, ZN 
                           => N3232);
   U16840 : OAI21_X1 port map( B1 => n1065_port, B2 => n11477, A => n11168, ZN 
                           => N3233);
   U16841 : OAI21_X1 port map( B1 => n1064_port, B2 => n11477, A => n11172, ZN 
                           => N3234);
   U16842 : OAI21_X1 port map( B1 => n1063_port, B2 => n11477, A => n11176, ZN 
                           => N3235);
   U16843 : OAI21_X1 port map( B1 => n1062_port, B2 => n11477, A => n11180, ZN 
                           => N3236);
   U16844 : OAI21_X1 port map( B1 => n1061_port, B2 => n11477, A => n11184, ZN 
                           => N3237);
   U16845 : OAI21_X1 port map( B1 => n1060_port, B2 => n11477, A => n11188, ZN 
                           => N3238);
   U16846 : OAI21_X1 port map( B1 => n1059_port, B2 => n11477, A => n11192, ZN 
                           => N3239);
   U16847 : OAI21_X1 port map( B1 => n1058_port, B2 => n11477, A => n11196, ZN 
                           => N3240);
   U16848 : OAI21_X1 port map( B1 => n1057_port, B2 => n11476, A => n11200, ZN 
                           => N3241);
   U16849 : OAI21_X1 port map( B1 => n1056_port, B2 => n11476, A => n11204, ZN 
                           => N3242);
   U16850 : OAI21_X1 port map( B1 => n1055_port, B2 => n11476, A => n11208, ZN 
                           => N3243);
   U16851 : OAI21_X1 port map( B1 => n1054_port, B2 => n11476, A => n11212, ZN 
                           => N3244);
   U16852 : OAI21_X1 port map( B1 => n1053_port, B2 => n11476, A => n11216, ZN 
                           => N3245);
   U16853 : OAI21_X1 port map( B1 => n1052_port, B2 => n11476, A => n11220, ZN 
                           => N3246);
   U16854 : OAI21_X1 port map( B1 => n1051_port, B2 => n11476, A => n11224, ZN 
                           => N3247);
   U16855 : OAI21_X1 port map( B1 => n1050_port, B2 => n11476, A => n11228, ZN 
                           => N3248);
   U16856 : OAI21_X1 port map( B1 => n1049_port, B2 => n11476, A => n11232, ZN 
                           => N3249);
   U16857 : OAI21_X1 port map( B1 => n1048_port, B2 => n11476, A => n11236, ZN 
                           => N3250);
   U16858 : OAI21_X1 port map( B1 => n1047_port, B2 => n11476, A => n11240, ZN 
                           => N3251);
   U16859 : OAI21_X1 port map( B1 => n1046_port, B2 => n11476, A => n11244, ZN 
                           => N3252);
   U16860 : OAI21_X1 port map( B1 => n1045_port, B2 => n11475, A => n11248, ZN 
                           => N3253);
   U16861 : OAI21_X1 port map( B1 => n1044_port, B2 => n11475, A => n11252, ZN 
                           => N3254);
   U16862 : OAI21_X1 port map( B1 => n1043_port, B2 => n11475, A => n11256, ZN 
                           => N3255);
   U16863 : OAI21_X1 port map( B1 => n1042_port, B2 => n11475, A => n11260, ZN 
                           => N3256);
   U16864 : OAI21_X1 port map( B1 => n1041_port, B2 => n11475, A => n11264, ZN 
                           => N3257);
   U16865 : OAI21_X1 port map( B1 => n1040_port, B2 => n11475, A => n11268, ZN 
                           => N3258);
   U16866 : OAI21_X1 port map( B1 => n1039_port, B2 => n11475, A => n11272, ZN 
                           => N3259);
   U16867 : OAI21_X1 port map( B1 => n1038_port, B2 => n11475, A => n11276, ZN 
                           => N3260);
   U16868 : OAI21_X1 port map( B1 => n1037_port, B2 => n11475, A => n11280, ZN 
                           => N3261);
   U16869 : OAI21_X1 port map( B1 => n1036_port, B2 => n11475, A => n11284, ZN 
                           => N3262);
   U16870 : OAI21_X1 port map( B1 => n1035_port, B2 => n11475, A => n11288, ZN 
                           => N3263);
   U16871 : OAI21_X1 port map( B1 => n1034_port, B2 => n11480, A => n11292, ZN 
                           => N3264);
   U16872 : OAI21_X1 port map( B1 => n1033_port, B2 => n11491, A => n11296, ZN 
                           => N3265);
   U16873 : OAI21_X1 port map( B1 => n1032_port, B2 => n11378, A => n11300, ZN 
                           => N3266);
   U16874 : OAI21_X1 port map( B1 => n1031_port, B2 => n11367, A => n11304, ZN 
                           => N3267);
   U16875 : OAI21_X1 port map( B1 => n1030_port, B2 => n11367, A => n11308, ZN 
                           => N3268);
   U16876 : OAI21_X1 port map( B1 => n1029_port, B2 => n11367, A => n11312, ZN 
                           => N3269);
   U16877 : OAI21_X1 port map( B1 => n1028_port, B2 => n11367, A => n11316, ZN 
                           => N3270);
   U16878 : OAI21_X1 port map( B1 => n1027_port, B2 => n11367, A => n11320, ZN 
                           => N3271);
   U16879 : OAI21_X1 port map( B1 => n1026_port, B2 => n11367, A => n11324, ZN 
                           => N3272);
   U16880 : OAI21_X1 port map( B1 => n1025_port, B2 => n11367, A => n11328, ZN 
                           => N3273);
   U16881 : OAI21_X1 port map( B1 => n1024_port, B2 => n11366, A => n11076, ZN 
                           => N3275);
   U16882 : OAI21_X1 port map( B1 => n1023_port, B2 => n11366, A => n11080, ZN 
                           => N3276);
   U16883 : OAI21_X1 port map( B1 => n1022_port, B2 => n11366, A => n11084, ZN 
                           => N3277);
   U16884 : OAI21_X1 port map( B1 => n1021_port, B2 => n11366, A => n11088, ZN 
                           => N3278);
   U16885 : OAI21_X1 port map( B1 => n1020_port, B2 => n11366, A => n11092, ZN 
                           => N3279);
   U16886 : OAI21_X1 port map( B1 => n1019_port, B2 => n11366, A => n11096, ZN 
                           => N3280);
   U16887 : OAI21_X1 port map( B1 => n1018_port, B2 => n11366, A => n11100, ZN 
                           => N3281);
   U16888 : OAI21_X1 port map( B1 => n1017_port, B2 => n11366, A => n11104, ZN 
                           => N3282);
   U16889 : OAI21_X1 port map( B1 => n1016_port, B2 => n11366, A => n11108, ZN 
                           => N3283);
   U16890 : OAI21_X1 port map( B1 => n1015_port, B2 => n11366, A => n11112, ZN 
                           => N3284);
   U16891 : OAI21_X1 port map( B1 => n1014_port, B2 => n11366, A => n11116, ZN 
                           => N3285);
   U16892 : OAI21_X1 port map( B1 => n1013_port, B2 => n11366, A => n11120, ZN 
                           => N3286);
   U16893 : OAI21_X1 port map( B1 => n1012_port, B2 => n11365, A => n11124, ZN 
                           => N3287);
   U16894 : OAI21_X1 port map( B1 => n1011_port, B2 => n11365, A => n11128, ZN 
                           => N3288);
   U16895 : OAI21_X1 port map( B1 => n1010_port, B2 => n11365, A => n11132, ZN 
                           => N3289);
   U16896 : OAI21_X1 port map( B1 => n1009_port, B2 => n11365, A => n11136, ZN 
                           => N3290);
   U16897 : OAI21_X1 port map( B1 => n1008_port, B2 => n11365, A => n11140, ZN 
                           => N3291);
   U16898 : OAI21_X1 port map( B1 => n1007_port, B2 => n11365, A => n11144, ZN 
                           => N3292);
   U16899 : OAI21_X1 port map( B1 => n1006_port, B2 => n11365, A => n11148, ZN 
                           => N3293);
   U16900 : OAI21_X1 port map( B1 => n1005_port, B2 => n11365, A => n11152, ZN 
                           => N3294);
   U16901 : OAI21_X1 port map( B1 => n1004_port, B2 => n11365, A => n11156, ZN 
                           => N3295);
   U16902 : OAI21_X1 port map( B1 => n1003_port, B2 => n11365, A => n11160, ZN 
                           => N3296);
   U16903 : OAI21_X1 port map( B1 => n1002_port, B2 => n11365, A => n11164, ZN 
                           => N3297);
   U16904 : OAI21_X1 port map( B1 => n1001_port, B2 => n11365, A => n11168, ZN 
                           => N3298);
   U16905 : OAI21_X1 port map( B1 => n1000_port, B2 => n11364, A => n11172, ZN 
                           => N3299);
   U16906 : OAI21_X1 port map( B1 => n999_port, B2 => n11364, A => n11176, ZN 
                           => N3300);
   U16907 : OAI21_X1 port map( B1 => n998_port, B2 => n11364, A => n11180, ZN 
                           => N3301);
   U16908 : OAI21_X1 port map( B1 => n997_port, B2 => n11364, A => n11184, ZN 
                           => N3302);
   U16909 : OAI21_X1 port map( B1 => n996_port, B2 => n11364, A => n11188, ZN 
                           => N3303);
   U16910 : OAI21_X1 port map( B1 => n995_port, B2 => n11364, A => n11192, ZN 
                           => N3304);
   U16911 : OAI21_X1 port map( B1 => n994_port, B2 => n11364, A => n11196, ZN 
                           => N3305);
   U16912 : OAI21_X1 port map( B1 => n993_port, B2 => n11364, A => n11200, ZN 
                           => N3306);
   U16913 : OAI21_X1 port map( B1 => n992_port, B2 => n11364, A => n11204, ZN 
                           => N3307);
   U16914 : OAI21_X1 port map( B1 => n991_port, B2 => n11364, A => n11208, ZN 
                           => N3308);
   U16915 : OAI21_X1 port map( B1 => n990_port, B2 => n11364, A => n11212, ZN 
                           => N3309);
   U16916 : OAI21_X1 port map( B1 => n989_port, B2 => n11364, A => n11216, ZN 
                           => N3310);
   U16917 : OAI21_X1 port map( B1 => n988_port, B2 => n11363, A => n11220, ZN 
                           => N3311);
   U16918 : OAI21_X1 port map( B1 => n987_port, B2 => n11363, A => n11224, ZN 
                           => N3312);
   U16919 : OAI21_X1 port map( B1 => n986_port, B2 => n11363, A => n11228, ZN 
                           => N3313);
   U16920 : OAI21_X1 port map( B1 => n985_port, B2 => n11363, A => n11232, ZN 
                           => N3314);
   U16921 : OAI21_X1 port map( B1 => n984_port, B2 => n11363, A => n11236, ZN 
                           => N3315);
   U16922 : OAI21_X1 port map( B1 => n983_port, B2 => n11363, A => n11240, ZN 
                           => N3316);
   U16923 : OAI21_X1 port map( B1 => n982_port, B2 => n11363, A => n11244, ZN 
                           => N3317);
   U16924 : OAI21_X1 port map( B1 => n981_port, B2 => n11363, A => n11248, ZN 
                           => N3318);
   U16925 : OAI21_X1 port map( B1 => n980_port, B2 => n11363, A => n11252, ZN 
                           => N3319);
   U16926 : OAI21_X1 port map( B1 => n979_port, B2 => n11363, A => n11256, ZN 
                           => N3320);
   U16927 : OAI21_X1 port map( B1 => n978_port, B2 => n11363, A => n11260, ZN 
                           => N3321);
   U16928 : OAI21_X1 port map( B1 => n977_port, B2 => n11363, A => n11264, ZN 
                           => N3322);
   U16929 : OAI21_X1 port map( B1 => n976_port, B2 => n11362, A => n11268, ZN 
                           => N3323);
   U16930 : OAI21_X1 port map( B1 => n975_port, B2 => n11362, A => n11272, ZN 
                           => N3324);
   U16931 : OAI21_X1 port map( B1 => n974_port, B2 => n11362, A => n11276, ZN 
                           => N3325);
   U16932 : OAI21_X1 port map( B1 => n973_port, B2 => n11362, A => n11280, ZN 
                           => N3326);
   U16933 : OAI21_X1 port map( B1 => n972_port, B2 => n11362, A => n11284, ZN 
                           => N3327);
   U16934 : OAI21_X1 port map( B1 => n971_port, B2 => n11362, A => n11288, ZN 
                           => N3328);
   U16935 : OAI21_X1 port map( B1 => n970_port, B2 => n11362, A => n11292, ZN 
                           => N3329);
   U16936 : OAI21_X1 port map( B1 => n969_port, B2 => n11362, A => n11296, ZN 
                           => N3330);
   U16937 : OAI21_X1 port map( B1 => n968_port, B2 => n11362, A => n11300, ZN 
                           => N3331);
   U16938 : OAI21_X1 port map( B1 => n967_port, B2 => n11362, A => n11304, ZN 
                           => N3332);
   U16939 : OAI21_X1 port map( B1 => n966_port, B2 => n11362, A => n11308, ZN 
                           => N3333);
   U16940 : OAI21_X1 port map( B1 => n965_port, B2 => n11361, A => n11312, ZN 
                           => N3334);
   U16941 : OAI21_X1 port map( B1 => n964_port, B2 => n11361, A => n11316, ZN 
                           => N3335);
   U16942 : OAI21_X1 port map( B1 => n963_port, B2 => n11361, A => n11320, ZN 
                           => N3336);
   U16943 : OAI21_X1 port map( B1 => n962_port, B2 => n11361, A => n11324, ZN 
                           => N3337);
   U16944 : OAI21_X1 port map( B1 => n961_port, B2 => n11361, A => n11328, ZN 
                           => N3338);
   U16945 : OAI21_X1 port map( B1 => n960_port, B2 => n11361, A => n11076, ZN 
                           => N3340);
   U16946 : OAI21_X1 port map( B1 => n959_port, B2 => n11361, A => n11080, ZN 
                           => N3341);
   U16947 : OAI21_X1 port map( B1 => n958_port, B2 => n11361, A => n11084, ZN 
                           => N3342);
   U16948 : OAI21_X1 port map( B1 => n957_port, B2 => n11361, A => n11088, ZN 
                           => N3343);
   U16949 : OAI21_X1 port map( B1 => n956_port, B2 => n11361, A => n11092, ZN 
                           => N3344);
   U16950 : OAI21_X1 port map( B1 => n955_port, B2 => n11361, A => n11096, ZN 
                           => N3345);
   U16951 : OAI21_X1 port map( B1 => n954_port, B2 => n11361, A => n11100, ZN 
                           => N3346);
   U16952 : OAI21_X1 port map( B1 => n953_port, B2 => n11360, A => n11104, ZN 
                           => N3347);
   U16953 : OAI21_X1 port map( B1 => n952_port, B2 => n11360, A => n11108, ZN 
                           => N3348);
   U16954 : OAI21_X1 port map( B1 => n951_port, B2 => n11360, A => n11112, ZN 
                           => N3349);
   U16955 : OAI21_X1 port map( B1 => n950_port, B2 => n11360, A => n11116, ZN 
                           => N3350);
   U16956 : OAI21_X1 port map( B1 => n949_port, B2 => n11360, A => n11120, ZN 
                           => N3351);
   U16957 : OAI21_X1 port map( B1 => n948_port, B2 => n11360, A => n11124, ZN 
                           => N3352);
   U16958 : OAI21_X1 port map( B1 => n947_port, B2 => n11360, A => n11128, ZN 
                           => N3353);
   U16959 : OAI21_X1 port map( B1 => n946_port, B2 => n11360, A => n11132, ZN 
                           => N3354);
   U16960 : OAI21_X1 port map( B1 => n945_port, B2 => n11360, A => n11136, ZN 
                           => N3355);
   U16961 : OAI21_X1 port map( B1 => n944_port, B2 => n11360, A => n11140, ZN 
                           => N3356);
   U16962 : OAI21_X1 port map( B1 => n943_port, B2 => n11360, A => n11144, ZN 
                           => N3357);
   U16963 : OAI21_X1 port map( B1 => n942_port, B2 => n11360, A => n11148, ZN 
                           => N3358);
   U16964 : OAI21_X1 port map( B1 => n941_port, B2 => n11359, A => n11152, ZN 
                           => N3359);
   U16965 : OAI21_X1 port map( B1 => n940_port, B2 => n11359, A => n11156, ZN 
                           => N3360);
   U16966 : OAI21_X1 port map( B1 => n939_port, B2 => n11359, A => n11160, ZN 
                           => N3361);
   U16967 : OAI21_X1 port map( B1 => n938_port, B2 => n11359, A => n11164, ZN 
                           => N3362);
   U16968 : OAI21_X1 port map( B1 => n937_port, B2 => n11359, A => n11168, ZN 
                           => N3363);
   U16969 : OAI21_X1 port map( B1 => n936_port, B2 => n11359, A => n11172, ZN 
                           => N3364);
   U16970 : OAI21_X1 port map( B1 => n935_port, B2 => n11359, A => n11176, ZN 
                           => N3365);
   U16971 : OAI21_X1 port map( B1 => n934_port, B2 => n11359, A => n11180, ZN 
                           => N3366);
   U16972 : OAI21_X1 port map( B1 => n933_port, B2 => n11359, A => n11184, ZN 
                           => N3367);
   U16973 : OAI21_X1 port map( B1 => n932_port, B2 => n11359, A => n11188, ZN 
                           => N3368);
   U16974 : OAI21_X1 port map( B1 => n931_port, B2 => n11359, A => n11192, ZN 
                           => N3369);
   U16975 : OAI21_X1 port map( B1 => n930_port, B2 => n11359, A => n11196, ZN 
                           => N3370);
   U16976 : OAI21_X1 port map( B1 => n929_port, B2 => n11358, A => n11200, ZN 
                           => N3371);
   U16977 : OAI21_X1 port map( B1 => n928_port, B2 => n11358, A => n11204, ZN 
                           => N3372);
   U16978 : OAI21_X1 port map( B1 => n927_port, B2 => n11358, A => n11208, ZN 
                           => N3373);
   U16979 : OAI21_X1 port map( B1 => n926_port, B2 => n11358, A => n11212, ZN 
                           => N3374);
   U16980 : OAI21_X1 port map( B1 => n925_port, B2 => n11358, A => n11216, ZN 
                           => N3375);
   U16981 : OAI21_X1 port map( B1 => n924_port, B2 => n11358, A => n11220, ZN 
                           => N3376);
   U16982 : OAI21_X1 port map( B1 => n923_port, B2 => n11358, A => n11224, ZN 
                           => N3377);
   U16983 : OAI21_X1 port map( B1 => n922_port, B2 => n11358, A => n11228, ZN 
                           => N3378);
   U16984 : OAI21_X1 port map( B1 => n921_port, B2 => n11358, A => n11232, ZN 
                           => N3379);
   U16985 : OAI21_X1 port map( B1 => n920_port, B2 => n11358, A => n11236, ZN 
                           => N3380);
   U16986 : OAI21_X1 port map( B1 => n919_port, B2 => n11358, A => n11240, ZN 
                           => N3381);
   U16987 : OAI21_X1 port map( B1 => n918_port, B2 => n11358, A => n11244, ZN 
                           => N3382);
   U16988 : OAI21_X1 port map( B1 => n917_port, B2 => n11357, A => n11248, ZN 
                           => N3383);
   U16989 : OAI21_X1 port map( B1 => n916_port, B2 => n11357, A => n11252, ZN 
                           => N3384);
   U16990 : OAI21_X1 port map( B1 => n915_port, B2 => n11357, A => n11256, ZN 
                           => N3385);
   U16991 : OAI21_X1 port map( B1 => n914_port, B2 => n11357, A => n11260, ZN 
                           => N3386);
   U16992 : OAI21_X1 port map( B1 => n913_port, B2 => n11357, A => n11264, ZN 
                           => N3387);
   U16993 : OAI21_X1 port map( B1 => n912_port, B2 => n11357, A => n11268, ZN 
                           => N3388);
   U16994 : OAI21_X1 port map( B1 => n911_port, B2 => n11357, A => n11272, ZN 
                           => N3389);
   U16995 : OAI21_X1 port map( B1 => n910_port, B2 => n11357, A => n11276, ZN 
                           => N3390);
   U16996 : OAI21_X1 port map( B1 => n909_port, B2 => n11357, A => n11280, ZN 
                           => N3391);
   U16997 : OAI21_X1 port map( B1 => n908_port, B2 => n11357, A => n11284, ZN 
                           => N3392);
   U16998 : OAI21_X1 port map( B1 => n907_port, B2 => n11357, A => n11288, ZN 
                           => N3393);
   U16999 : OAI21_X1 port map( B1 => n906_port, B2 => n11357, A => n11292, ZN 
                           => N3394);
   U17000 : OAI21_X1 port map( B1 => n905_port, B2 => n11356, A => n11296, ZN 
                           => N3395);
   U17001 : OAI21_X1 port map( B1 => n904_port, B2 => n11356, A => n11300, ZN 
                           => N3396);
   U17002 : OAI21_X1 port map( B1 => n903_port, B2 => n11362, A => n11304, ZN 
                           => N3397);
   U17003 : OAI21_X1 port map( B1 => n902_port, B2 => n11378, A => n11308, ZN 
                           => N3398);
   U17004 : OAI21_X1 port map( B1 => n901_port, B2 => n11378, A => n11312, ZN 
                           => N3399);
   U17005 : OAI21_X1 port map( B1 => n900_port, B2 => n11378, A => n11316, ZN 
                           => N3400);
   U17006 : OAI21_X1 port map( B1 => n899_port, B2 => n11377, A => n11320, ZN 
                           => N3401);
   U17007 : OAI21_X1 port map( B1 => n898_port, B2 => n11377, A => n11324, ZN 
                           => N3402);
   U17008 : OAI21_X1 port map( B1 => n897_port, B2 => n11377, A => n11328, ZN 
                           => N3403);
   U17009 : OAI21_X1 port map( B1 => n896_port, B2 => n11377, A => n11076, ZN 
                           => N3405);
   U17010 : OAI21_X1 port map( B1 => n895_port, B2 => n11377, A => n11080, ZN 
                           => N3406);
   U17011 : OAI21_X1 port map( B1 => n894_port, B2 => n11377, A => n11084, ZN 
                           => N3407);
   U17012 : OAI21_X1 port map( B1 => n893_port, B2 => n11377, A => n11088, ZN 
                           => N3408);
   U17013 : OAI21_X1 port map( B1 => n892_port, B2 => n11377, A => n11092, ZN 
                           => N3409);
   U17014 : OAI21_X1 port map( B1 => n891_port, B2 => n11377, A => n11096, ZN 
                           => N3410);
   U17015 : OAI21_X1 port map( B1 => n890_port, B2 => n11377, A => n11100, ZN 
                           => N3411);
   U17016 : OAI21_X1 port map( B1 => n889_port, B2 => n11377, A => n11104, ZN 
                           => N3412);
   U17017 : OAI21_X1 port map( B1 => n888_port, B2 => n11377, A => n11108, ZN 
                           => N3413);
   U17018 : OAI21_X1 port map( B1 => n887_port, B2 => n11376, A => n11112, ZN 
                           => N3414);
   U17019 : OAI21_X1 port map( B1 => n886_port, B2 => n11376, A => n11116, ZN 
                           => N3415);
   U17020 : OAI21_X1 port map( B1 => n885_port, B2 => n11376, A => n11120, ZN 
                           => N3416);
   U17021 : OAI21_X1 port map( B1 => n884_port, B2 => n11376, A => n11124, ZN 
                           => N3417);
   U17022 : OAI21_X1 port map( B1 => n883_port, B2 => n11376, A => n11128, ZN 
                           => N3418);
   U17023 : OAI21_X1 port map( B1 => n882_port, B2 => n11376, A => n11132, ZN 
                           => N3419);
   U17024 : OAI21_X1 port map( B1 => n881_port, B2 => n11376, A => n11136, ZN 
                           => N3420);
   U17025 : OAI21_X1 port map( B1 => n880_port, B2 => n11376, A => n11140, ZN 
                           => N3421);
   U17026 : OAI21_X1 port map( B1 => n879_port, B2 => n11376, A => n11144, ZN 
                           => N3422);
   U17027 : OAI21_X1 port map( B1 => n878_port, B2 => n11376, A => n11148, ZN 
                           => N3423);
   U17028 : OAI21_X1 port map( B1 => n877_port, B2 => n11376, A => n11152, ZN 
                           => N3424);
   U17029 : OAI21_X1 port map( B1 => n876_port, B2 => n11376, A => n11156, ZN 
                           => N3425);
   U17030 : OAI21_X1 port map( B1 => n875_port, B2 => n11375, A => n11160, ZN 
                           => N3426);
   U17031 : OAI21_X1 port map( B1 => n874_port, B2 => n11375, A => n11164, ZN 
                           => N3427);
   U17032 : OAI21_X1 port map( B1 => n873_port, B2 => n11375, A => n11168, ZN 
                           => N3428);
   U17033 : OAI21_X1 port map( B1 => n872_port, B2 => n11375, A => n11172, ZN 
                           => N3429);
   U17034 : OAI21_X1 port map( B1 => n871_port, B2 => n11375, A => n11176, ZN 
                           => N3430);
   U17035 : OAI21_X1 port map( B1 => n870_port, B2 => n11375, A => n11180, ZN 
                           => N3431);
   U17036 : OAI21_X1 port map( B1 => n869_port, B2 => n11375, A => n11184, ZN 
                           => N3432);
   U17037 : OAI21_X1 port map( B1 => n868_port, B2 => n11375, A => n11188, ZN 
                           => N3433);
   U17038 : OAI21_X1 port map( B1 => n867_port, B2 => n11375, A => n11192, ZN 
                           => N3434);
   U17039 : OAI21_X1 port map( B1 => n866_port, B2 => n11375, A => n11196, ZN 
                           => N3435);
   U17040 : OAI21_X1 port map( B1 => n865_port, B2 => n11375, A => n11200, ZN 
                           => N3436);
   U17041 : OAI21_X1 port map( B1 => n864_port, B2 => n11375, A => n11204, ZN 
                           => N3437);
   U17042 : OAI21_X1 port map( B1 => n863_port, B2 => n11374, A => n11208, ZN 
                           => N3438);
   U17043 : OAI21_X1 port map( B1 => n862_port, B2 => n11374, A => n11212, ZN 
                           => N3439);
   U17044 : OAI21_X1 port map( B1 => n861_port, B2 => n11374, A => n11216, ZN 
                           => N3440);
   U17045 : OAI21_X1 port map( B1 => n860_port, B2 => n11374, A => n11220, ZN 
                           => N3441);
   U17046 : OAI21_X1 port map( B1 => n859_port, B2 => n11374, A => n11224, ZN 
                           => N3442);
   U17047 : OAI21_X1 port map( B1 => n858_port, B2 => n11374, A => n11228, ZN 
                           => N3443);
   U17048 : OAI21_X1 port map( B1 => n857_port, B2 => n11374, A => n11232, ZN 
                           => N3444);
   U17049 : OAI21_X1 port map( B1 => n856_port, B2 => n11374, A => n11236, ZN 
                           => N3445);
   U17050 : OAI21_X1 port map( B1 => n855_port, B2 => n11374, A => n11240, ZN 
                           => N3446);
   U17051 : OAI21_X1 port map( B1 => n854_port, B2 => n11374, A => n11244, ZN 
                           => N3447);
   U17052 : OAI21_X1 port map( B1 => n853_port, B2 => n11374, A => n11248, ZN 
                           => N3448);
   U17053 : OAI21_X1 port map( B1 => n852_port, B2 => n11374, A => n11252, ZN 
                           => N3449);
   U17054 : OAI21_X1 port map( B1 => n851_port, B2 => n11373, A => n11256, ZN 
                           => N3450);
   U17055 : OAI21_X1 port map( B1 => n850_port, B2 => n11373, A => n11260, ZN 
                           => N3451);
   U17056 : OAI21_X1 port map( B1 => n849_port, B2 => n11373, A => n11264, ZN 
                           => N3452);
   U17057 : OAI21_X1 port map( B1 => n848_port, B2 => n11373, A => n11268, ZN 
                           => N3453);
   U17058 : OAI21_X1 port map( B1 => n847_port, B2 => n11373, A => n11272, ZN 
                           => N3454);
   U17059 : OAI21_X1 port map( B1 => n846_port, B2 => n11373, A => n11276, ZN 
                           => N3455);
   U17060 : OAI21_X1 port map( B1 => n845_port, B2 => n11373, A => n11280, ZN 
                           => N3456);
   U17061 : OAI21_X1 port map( B1 => n844_port, B2 => n11373, A => n11284, ZN 
                           => N3457);
   U17062 : OAI21_X1 port map( B1 => n843_port, B2 => n11373, A => n11288, ZN 
                           => N3458);
   U17063 : OAI21_X1 port map( B1 => n842_port, B2 => n11373, A => n11292, ZN 
                           => N3459);
   U17064 : OAI21_X1 port map( B1 => n841_port, B2 => n11373, A => n11296, ZN 
                           => N3460);
   U17065 : OAI21_X1 port map( B1 => n840_port, B2 => n11373, A => n11300, ZN 
                           => N3461);
   U17066 : OAI21_X1 port map( B1 => n839_port, B2 => n11372, A => n11304, ZN 
                           => N3462);
   U17067 : OAI21_X1 port map( B1 => n838_port, B2 => n11372, A => n11308, ZN 
                           => N3463);
   U17068 : OAI21_X1 port map( B1 => n837_port, B2 => n11372, A => n11312, ZN 
                           => N3464);
   U17069 : OAI21_X1 port map( B1 => n836_port, B2 => n11372, A => n11316, ZN 
                           => N3465);
   U17070 : OAI21_X1 port map( B1 => n835_port, B2 => n11372, A => n11320, ZN 
                           => N3466);
   U17071 : OAI21_X1 port map( B1 => n834_port, B2 => n11372, A => n11324, ZN 
                           => N3467);
   U17072 : OAI21_X1 port map( B1 => n833_port, B2 => n11372, A => n11328, ZN 
                           => N3468);
   U17073 : OAI21_X1 port map( B1 => n832_port, B2 => n11372, A => n11076, ZN 
                           => N3470);
   U17074 : OAI21_X1 port map( B1 => n831_port, B2 => n11372, A => n11080, ZN 
                           => N3471);
   U17075 : OAI21_X1 port map( B1 => n830_port, B2 => n11372, A => n11084, ZN 
                           => N3472);
   U17076 : OAI21_X1 port map( B1 => n829_port, B2 => n11372, A => n11088, ZN 
                           => N3473);
   U17077 : OAI21_X1 port map( B1 => n828_port, B2 => n11371, A => n11092, ZN 
                           => N3474);
   U17078 : OAI21_X1 port map( B1 => n827_port, B2 => n11371, A => n11096, ZN 
                           => N3475);
   U17079 : OAI21_X1 port map( B1 => n826_port, B2 => n11371, A => n11100, ZN 
                           => N3476);
   U17080 : OAI21_X1 port map( B1 => n825_port, B2 => n11371, A => n11104, ZN 
                           => N3477);
   U17081 : OAI21_X1 port map( B1 => n824_port, B2 => n11371, A => n11108, ZN 
                           => N3478);
   U17082 : OAI21_X1 port map( B1 => n823_port, B2 => n11371, A => n11112, ZN 
                           => N3479);
   U17083 : OAI21_X1 port map( B1 => n822_port, B2 => n11371, A => n11116, ZN 
                           => N3480);
   U17084 : OAI21_X1 port map( B1 => n821_port, B2 => n11371, A => n11120, ZN 
                           => N3481);
   U17085 : OAI21_X1 port map( B1 => n820_port, B2 => n11371, A => n11124, ZN 
                           => N3482);
   U17086 : OAI21_X1 port map( B1 => n819_port, B2 => n11371, A => n11128, ZN 
                           => N3483);
   U17087 : OAI21_X1 port map( B1 => n818_port, B2 => n11371, A => n11132, ZN 
                           => N3484);
   U17088 : OAI21_X1 port map( B1 => n817_port, B2 => n11371, A => n11136, ZN 
                           => N3485);
   U17089 : OAI21_X1 port map( B1 => n816_port, B2 => n11370, A => n11140, ZN 
                           => N3486);
   U17090 : OAI21_X1 port map( B1 => n815_port, B2 => n11370, A => n11144, ZN 
                           => N3487);
   U17091 : OAI21_X1 port map( B1 => n814_port, B2 => n11370, A => n11148, ZN 
                           => N3488);
   U17092 : OAI21_X1 port map( B1 => n813_port, B2 => n11370, A => n11152, ZN 
                           => N3489);
   U17093 : OAI21_X1 port map( B1 => n812_port, B2 => n11370, A => n11156, ZN 
                           => N3490);
   U17094 : OAI21_X1 port map( B1 => n811_port, B2 => n11370, A => n11160, ZN 
                           => N3491);
   U17095 : OAI21_X1 port map( B1 => n810_port, B2 => n11370, A => n11164, ZN 
                           => N3492);
   U17096 : OAI21_X1 port map( B1 => n809_port, B2 => n11370, A => n11168, ZN 
                           => N3493);
   U17097 : OAI21_X1 port map( B1 => n808_port, B2 => n11370, A => n11172, ZN 
                           => N3494);
   U17098 : OAI21_X1 port map( B1 => n807_port, B2 => n11370, A => n11176, ZN 
                           => N3495);
   U17099 : OAI21_X1 port map( B1 => n806_port, B2 => n11370, A => n11180, ZN 
                           => N3496);
   U17100 : OAI21_X1 port map( B1 => n805_port, B2 => n11370, A => n11184, ZN 
                           => N3497);
   U17101 : OAI21_X1 port map( B1 => n804_port, B2 => n11369, A => n11188, ZN 
                           => N3498);
   U17102 : OAI21_X1 port map( B1 => n803_port, B2 => n11369, A => n11192, ZN 
                           => N3499);
   U17103 : OAI21_X1 port map( B1 => n802_port, B2 => n11369, A => n11196, ZN 
                           => N3500);
   U17104 : OAI21_X1 port map( B1 => n801_port, B2 => n11369, A => n11200, ZN 
                           => N3501);
   U17105 : OAI21_X1 port map( B1 => n800_port, B2 => n11369, A => n11204, ZN 
                           => N3502);
   U17106 : OAI21_X1 port map( B1 => n799_port, B2 => n11369, A => n11208, ZN 
                           => N3503);
   U17107 : OAI21_X1 port map( B1 => n798_port, B2 => n11369, A => n11212, ZN 
                           => N3504);
   U17108 : OAI21_X1 port map( B1 => n797_port, B2 => n11369, A => n11216, ZN 
                           => N3505);
   U17109 : OAI21_X1 port map( B1 => n796_port, B2 => n11369, A => n11220, ZN 
                           => N3506);
   U17110 : OAI21_X1 port map( B1 => n795_port, B2 => n11369, A => n11224, ZN 
                           => N3507);
   U17111 : OAI21_X1 port map( B1 => n794_port, B2 => n11369, A => n11228, ZN 
                           => N3508);
   U17112 : OAI21_X1 port map( B1 => n793_port, B2 => n11369, A => n11232, ZN 
                           => N3509);
   U17113 : OAI21_X1 port map( B1 => n792_port, B2 => n11368, A => n11236, ZN 
                           => N3510);
   U17114 : OAI21_X1 port map( B1 => n791_port, B2 => n11368, A => n11240, ZN 
                           => N3511);
   U17115 : OAI21_X1 port map( B1 => n790_port, B2 => n11368, A => n11244, ZN 
                           => N3512);
   U17116 : OAI21_X1 port map( B1 => n789_port, B2 => n11368, A => n11248, ZN 
                           => N3513);
   U17117 : OAI21_X1 port map( B1 => n788_port, B2 => n11368, A => n11252, ZN 
                           => N3514);
   U17118 : OAI21_X1 port map( B1 => n787_port, B2 => n11368, A => n11256, ZN 
                           => N3515);
   U17119 : OAI21_X1 port map( B1 => n786_port, B2 => n11368, A => n11260, ZN 
                           => N3516);
   U17120 : OAI21_X1 port map( B1 => n785_port, B2 => n11368, A => n11264, ZN 
                           => N3517);
   U17121 : OAI21_X1 port map( B1 => n784_port, B2 => n11368, A => n11268, ZN 
                           => N3518);
   U17122 : OAI21_X1 port map( B1 => n783_port, B2 => n11368, A => n11272, ZN 
                           => N3519);
   U17123 : OAI21_X1 port map( B1 => n782_port, B2 => n11368, A => n11276, ZN 
                           => N3520);
   U17124 : OAI21_X1 port map( B1 => n781_port, B2 => n11368, A => n11280, ZN 
                           => N3521);
   U17125 : OAI21_X1 port map( B1 => n780_port, B2 => n11367, A => n11284, ZN 
                           => N3522);
   U17126 : OAI21_X1 port map( B1 => n779_port, B2 => n11367, A => n11288, ZN 
                           => N3523);
   U17127 : OAI21_X1 port map( B1 => n778_port, B2 => n11367, A => n11292, ZN 
                           => N3524);
   U17128 : OAI21_X1 port map( B1 => n777_port, B2 => n11367, A => n11296, ZN 
                           => N3525);
   U17129 : OAI21_X1 port map( B1 => n776_port, B2 => n11367, A => n11300, ZN 
                           => N3526);
   U17130 : OAI21_X1 port map( B1 => n775_port, B2 => n11372, A => n11304, ZN 
                           => N3527);
   U17131 : OAI21_X1 port map( B1 => n774_port, B2 => n11346, A => n11308, ZN 
                           => N3528);
   U17132 : OAI21_X1 port map( B1 => n773_port, B2 => n11345, A => n11312, ZN 
                           => N3529);
   U17133 : OAI21_X1 port map( B1 => n772_port, B2 => n11345, A => n11316, ZN 
                           => N3530);
   U17134 : OAI21_X1 port map( B1 => n771_port, B2 => n11345, A => n11320, ZN 
                           => N3531);
   U17135 : OAI21_X1 port map( B1 => n770_port, B2 => n11345, A => n11324, ZN 
                           => N3532);
   U17136 : OAI21_X1 port map( B1 => n769_port, B2 => n11345, A => n11328, ZN 
                           => N3533);
   U17137 : OAI21_X1 port map( B1 => n768_port, B2 => n11345, A => n11076, ZN 
                           => N3535);
   U17138 : OAI21_X1 port map( B1 => n767_port, B2 => n11345, A => n11080, ZN 
                           => N3536);
   U17139 : OAI21_X1 port map( B1 => n766_port, B2 => n11345, A => n11084, ZN 
                           => N3537);
   U17140 : OAI21_X1 port map( B1 => n765_port, B2 => n11345, A => n11088, ZN 
                           => N3538);
   U17141 : OAI21_X1 port map( B1 => n764_port, B2 => n11345, A => n11092, ZN 
                           => N3539);
   U17142 : OAI21_X1 port map( B1 => n763_port, B2 => n11345, A => n11096, ZN 
                           => N3540);
   U17143 : OAI21_X1 port map( B1 => n762_port, B2 => n11345, A => n11100, ZN 
                           => N3541);
   U17144 : OAI21_X1 port map( B1 => n761_port, B2 => n11344, A => n11104, ZN 
                           => N3542);
   U17145 : OAI21_X1 port map( B1 => n760_port, B2 => n11344, A => n11108, ZN 
                           => N3543);
   U17146 : OAI21_X1 port map( B1 => n759_port, B2 => n11344, A => n11112, ZN 
                           => N3544);
   U17147 : OAI21_X1 port map( B1 => n758_port, B2 => n11344, A => n11116, ZN 
                           => N3545);
   U17148 : OAI21_X1 port map( B1 => n757_port, B2 => n11344, A => n11120, ZN 
                           => N3546);
   U17149 : OAI21_X1 port map( B1 => n756_port, B2 => n11344, A => n11124, ZN 
                           => N3547);
   U17150 : OAI21_X1 port map( B1 => n755_port, B2 => n11344, A => n11128, ZN 
                           => N3548);
   U17151 : OAI21_X1 port map( B1 => n754_port, B2 => n11344, A => n11132, ZN 
                           => N3549);
   U17152 : OAI21_X1 port map( B1 => n753_port, B2 => n11344, A => n11136, ZN 
                           => N3550);
   U17153 : OAI21_X1 port map( B1 => n752_port, B2 => n11344, A => n11140, ZN 
                           => N3551);
   U17154 : OAI21_X1 port map( B1 => n751_port, B2 => n11344, A => n11144, ZN 
                           => N3552);
   U17155 : OAI21_X1 port map( B1 => n750_port, B2 => n11344, A => n11148, ZN 
                           => N3553);
   U17156 : OAI21_X1 port map( B1 => n749_port, B2 => n11343, A => n11152, ZN 
                           => N3554);
   U17157 : OAI21_X1 port map( B1 => n748_port, B2 => n11343, A => n11156, ZN 
                           => N3555);
   U17158 : OAI21_X1 port map( B1 => n747_port, B2 => n11343, A => n11160, ZN 
                           => N3556);
   U17159 : OAI21_X1 port map( B1 => n746_port, B2 => n11343, A => n11164, ZN 
                           => N3557);
   U17160 : OAI21_X1 port map( B1 => n745_port, B2 => n11343, A => n11168, ZN 
                           => N3558);
   U17161 : OAI21_X1 port map( B1 => n744_port, B2 => n11343, A => n11172, ZN 
                           => N3559);
   U17162 : OAI21_X1 port map( B1 => n743_port, B2 => n11343, A => n11176, ZN 
                           => N3560);
   U17163 : OAI21_X1 port map( B1 => n742_port, B2 => n11343, A => n11180, ZN 
                           => N3561);
   U17164 : OAI21_X1 port map( B1 => n741_port, B2 => n11343, A => n11184, ZN 
                           => N3562);
   U17165 : OAI21_X1 port map( B1 => n740_port, B2 => n11343, A => n11188, ZN 
                           => N3563);
   U17166 : OAI21_X1 port map( B1 => n739_port, B2 => n11343, A => n11192, ZN 
                           => N3564);
   U17167 : OAI21_X1 port map( B1 => n738_port, B2 => n11343, A => n11196, ZN 
                           => N3565);
   U17168 : OAI21_X1 port map( B1 => n737_port, B2 => n11342, A => n11200, ZN 
                           => N3566);
   U17169 : OAI21_X1 port map( B1 => n736_port, B2 => n11342, A => n11204, ZN 
                           => N3567);
   U17170 : OAI21_X1 port map( B1 => n735_port, B2 => n11342, A => n11208, ZN 
                           => N3568);
   U17171 : OAI21_X1 port map( B1 => n734_port, B2 => n11342, A => n11212, ZN 
                           => N3569);
   U17172 : OAI21_X1 port map( B1 => n733_port, B2 => n11342, A => n11216, ZN 
                           => N3570);
   U17173 : OAI21_X1 port map( B1 => n732_port, B2 => n11342, A => n11220, ZN 
                           => N3571);
   U17174 : OAI21_X1 port map( B1 => n731_port, B2 => n11342, A => n11224, ZN 
                           => N3572);
   U17175 : OAI21_X1 port map( B1 => n730_port, B2 => n11342, A => n11228, ZN 
                           => N3573);
   U17176 : OAI21_X1 port map( B1 => n729_port, B2 => n11342, A => n11232, ZN 
                           => N3574);
   U17177 : OAI21_X1 port map( B1 => n728_port, B2 => n11342, A => n11236, ZN 
                           => N3575);
   U17178 : OAI21_X1 port map( B1 => n727_port, B2 => n11342, A => n11240, ZN 
                           => N3576);
   U17179 : OAI21_X1 port map( B1 => n726_port, B2 => n11342, A => n11244, ZN 
                           => N3577);
   U17180 : OAI21_X1 port map( B1 => n725_port, B2 => n11341, A => n11248, ZN 
                           => N3578);
   U17181 : OAI21_X1 port map( B1 => n724_port, B2 => n11341, A => n11252, ZN 
                           => N3579);
   U17182 : OAI21_X1 port map( B1 => n723_port, B2 => n11341, A => n11256, ZN 
                           => N3580);
   U17183 : OAI21_X1 port map( B1 => n722_port, B2 => n11341, A => n11260, ZN 
                           => N3581);
   U17184 : OAI21_X1 port map( B1 => n721_port, B2 => n11341, A => n11264, ZN 
                           => N3582);
   U17185 : OAI21_X1 port map( B1 => n720_port, B2 => n11341, A => n11268, ZN 
                           => N3583);
   U17186 : OAI21_X1 port map( B1 => n719_port, B2 => n11341, A => n11272, ZN 
                           => N3584);
   U17187 : OAI21_X1 port map( B1 => n718_port, B2 => n11341, A => n11276, ZN 
                           => N3585);
   U17188 : OAI21_X1 port map( B1 => n717_port, B2 => n11341, A => n11280, ZN 
                           => N3586);
   U17189 : OAI21_X1 port map( B1 => n716_port, B2 => n11341, A => n11284, ZN 
                           => N3587);
   U17190 : OAI21_X1 port map( B1 => n715_port, B2 => n11341, A => n11288, ZN 
                           => N3588);
   U17191 : OAI21_X1 port map( B1 => n714_port, B2 => n11341, A => n11292, ZN 
                           => N3589);
   U17192 : OAI21_X1 port map( B1 => n713_port, B2 => n11340, A => n11296, ZN 
                           => N3590);
   U17193 : OAI21_X1 port map( B1 => n712_port, B2 => n11340, A => n11300, ZN 
                           => N3591);
   U17194 : OAI21_X1 port map( B1 => n711_port, B2 => n11340, A => n11304, ZN 
                           => N3592);
   U17195 : OAI21_X1 port map( B1 => n710_port, B2 => n11340, A => n11308, ZN 
                           => N3593);
   U17196 : OAI21_X1 port map( B1 => n709_port, B2 => n11340, A => n11312, ZN 
                           => N3594);
   U17197 : OAI21_X1 port map( B1 => n708_port, B2 => n11340, A => n11316, ZN 
                           => N3595);
   U17198 : OAI21_X1 port map( B1 => n707_port, B2 => n11340, A => n11320, ZN 
                           => N3596);
   U17199 : OAI21_X1 port map( B1 => n706_port, B2 => n11340, A => n11324, ZN 
                           => N3597);
   U17200 : OAI21_X1 port map( B1 => n705_port, B2 => n11339, A => n11328, ZN 
                           => N3598);
   U17201 : OAI21_X1 port map( B1 => n704_port, B2 => n11339, A => n11076, ZN 
                           => N3600);
   U17202 : OAI21_X1 port map( B1 => n703_port, B2 => n11339, A => n11080, ZN 
                           => N3601);
   U17203 : OAI21_X1 port map( B1 => n702_port, B2 => n11339, A => n11084, ZN 
                           => N3602);
   U17204 : OAI21_X1 port map( B1 => n701_port, B2 => n11339, A => n11088, ZN 
                           => N3603);
   U17205 : OAI21_X1 port map( B1 => n700_port, B2 => n11339, A => n11092, ZN 
                           => N3604);
   U17206 : OAI21_X1 port map( B1 => n699_port, B2 => n11338, A => n11096, ZN 
                           => N3605);
   U17207 : OAI21_X1 port map( B1 => n698_port, B2 => n11338, A => n11100, ZN 
                           => N3606);
   U17208 : OAI21_X1 port map( B1 => n697_port, B2 => n11339, A => n11104, ZN 
                           => N3607);
   U17209 : OAI21_X1 port map( B1 => n696_port, B2 => n11338, A => n11108, ZN 
                           => N3608);
   U17210 : OAI21_X1 port map( B1 => n695_port, B2 => n11338, A => n11112, ZN 
                           => N3609);
   U17211 : OAI21_X1 port map( B1 => n694_port, B2 => n11338, A => n11116, ZN 
                           => N3610);
   U17212 : OAI21_X1 port map( B1 => n693_port, B2 => n11338, A => n11120, ZN 
                           => N3611);
   U17213 : OAI21_X1 port map( B1 => n692_port, B2 => n11337, A => n11124, ZN 
                           => N3612);
   U17214 : OAI21_X1 port map( B1 => n691_port, B2 => n11338, A => n11128, ZN 
                           => N3613);
   U17215 : OAI21_X1 port map( B1 => n690_port, B2 => n11337, A => n11132, ZN 
                           => N3614);
   U17216 : OAI21_X1 port map( B1 => n689_port, B2 => n11337, A => n11136, ZN 
                           => N3615);
   U17217 : OAI21_X1 port map( B1 => n688_port, B2 => n11337, A => n11140, ZN 
                           => N3616);
   U17218 : OAI21_X1 port map( B1 => n687_port, B2 => n11337, A => n11144, ZN 
                           => N3617);
   U17219 : OAI21_X1 port map( B1 => n686_port, B2 => n11338, A => n11148, ZN 
                           => N3618);
   U17220 : OAI21_X1 port map( B1 => n685_port, B2 => n11338, A => n11152, ZN 
                           => N3619);
   U17221 : OAI21_X1 port map( B1 => n684_port, B2 => n11336, A => n11156, ZN 
                           => N3620);
   U17222 : OAI21_X1 port map( B1 => n683_port, B2 => n11336, A => n11160, ZN 
                           => N3621);
   U17223 : OAI21_X1 port map( B1 => n682_port, B2 => n11337, A => n11164, ZN 
                           => N3622);
   U17224 : OAI21_X1 port map( B1 => n681_port, B2 => n11336, A => n11168, ZN 
                           => N3623);
   U17225 : OAI21_X1 port map( B1 => n680_port, B2 => n11336, A => n11172, ZN 
                           => N3624);
   U17226 : OAI21_X1 port map( B1 => n679_port, B2 => n11336, A => n11176, ZN 
                           => N3625);
   U17227 : OAI21_X1 port map( B1 => n676_port, B2 => n11336, A => n11188, ZN 
                           => N3628);
   U17228 : OAI21_X1 port map( B1 => n673_port, B2 => n11336, A => n11200, ZN 
                           => N3631);
   U17229 : OAI21_X1 port map( B1 => n672_port, B2 => n11336, A => n11204, ZN 
                           => N3632);
   U17230 : OAI21_X1 port map( B1 => n670_port, B2 => n11336, A => n11212, ZN 
                           => N3634);
   U17231 : OAI21_X1 port map( B1 => n668_port, B2 => n11336, A => n11220, ZN 
                           => N3636);
   U17232 : OAI21_X1 port map( B1 => n666_port, B2 => n11337, A => n11228, ZN 
                           => N3638);
   U17233 : OAI21_X1 port map( B1 => n665_port, B2 => n11336, A => n11232, ZN 
                           => N3639);
   U17234 : OAI21_X1 port map( B1 => n664_port, B2 => n11337, A => n11236, ZN 
                           => N3640);
   U17235 : OAI21_X1 port map( B1 => n662_port, B2 => n11337, A => n11244, ZN 
                           => N3642);
   U17236 : OAI21_X1 port map( B1 => n661_port, B2 => n11338, A => n11248, ZN 
                           => N3643);
   U17237 : OAI21_X1 port map( B1 => n660_port, B2 => n11336, A => n11252, ZN 
                           => N3644);
   U17238 : OAI21_X1 port map( B1 => n659_port, B2 => n11337, A => n11256, ZN 
                           => N3645);
   U17239 : OAI21_X1 port map( B1 => n658_port, B2 => n11337, A => n11260, ZN 
                           => N3646);
   U17240 : OAI21_X1 port map( B1 => n657_port, B2 => n11337, A => n11264, ZN 
                           => N3647);
   U17241 : OAI21_X1 port map( B1 => n656_port, B2 => n11338, A => n11268, ZN 
                           => N3648);
   U17242 : OAI21_X1 port map( B1 => n655_port, B2 => n11338, A => n11272, ZN 
                           => N3649);
   U17243 : OAI21_X1 port map( B1 => n654_port, B2 => n11339, A => n11276, ZN 
                           => N3650);
   U17244 : OAI21_X1 port map( B1 => n653_port, B2 => n11339, A => n11280, ZN 
                           => N3651);
   U17245 : OAI21_X1 port map( B1 => n652_port, B2 => n11339, A => n11284, ZN 
                           => N3652);
   U17246 : OAI21_X1 port map( B1 => n651_port, B2 => n11339, A => n11288, ZN 
                           => N3653);
   U17247 : OAI21_X1 port map( B1 => n650_port, B2 => n11339, A => n11292, ZN 
                           => N3654);
   U17248 : OAI21_X1 port map( B1 => n649_port, B2 => n11340, A => n11296, ZN 
                           => N3655);
   U17249 : OAI21_X1 port map( B1 => n648_port, B2 => n11340, A => n11300, ZN 
                           => N3656);
   U17250 : OAI21_X1 port map( B1 => n647_port, B2 => n11340, A => n11304, ZN 
                           => N3657);
   U17251 : OAI21_X1 port map( B1 => n646_port, B2 => n11356, A => n11308, ZN 
                           => N3658);
   U17252 : OAI21_X1 port map( B1 => n645_port, B2 => n11356, A => n11312, ZN 
                           => N3659);
   U17253 : OAI21_X1 port map( B1 => n644_port, B2 => n11356, A => n11316, ZN 
                           => N3660);
   U17254 : OAI21_X1 port map( B1 => n643_port, B2 => n11356, A => n11320, ZN 
                           => N3661);
   U17255 : OAI21_X1 port map( B1 => n642_port, B2 => n11356, A => n11324, ZN 
                           => N3662);
   U17256 : OAI21_X1 port map( B1 => n641_port, B2 => n11356, A => n11328, ZN 
                           => N3663);
   U17257 : OAI21_X1 port map( B1 => n640_port, B2 => n11356, A => n11076, ZN 
                           => N3665);
   U17258 : OAI21_X1 port map( B1 => n639_port, B2 => n11356, A => n11080, ZN 
                           => N3666);
   U17259 : OAI21_X1 port map( B1 => n638_port, B2 => n11356, A => n11084, ZN 
                           => N3667);
   U17260 : OAI21_X1 port map( B1 => n637_port, B2 => n11355, A => n11088, ZN 
                           => N3668);
   U17261 : OAI21_X1 port map( B1 => n636_port, B2 => n11355, A => n11092, ZN 
                           => N3669);
   U17262 : OAI21_X1 port map( B1 => n635_port, B2 => n11355, A => n11096, ZN 
                           => N3670);
   U17263 : OAI21_X1 port map( B1 => n634_port, B2 => n11355, A => n11100, ZN 
                           => N3671);
   U17264 : OAI21_X1 port map( B1 => n633_port, B2 => n11355, A => n11104, ZN 
                           => N3672);
   U17265 : OAI21_X1 port map( B1 => n632_port, B2 => n11355, A => n11108, ZN 
                           => N3673);
   U17266 : OAI21_X1 port map( B1 => n631_port, B2 => n11355, A => n11112, ZN 
                           => N3674);
   U17267 : OAI21_X1 port map( B1 => n630_port, B2 => n11355, A => n11116, ZN 
                           => N3675);
   U17268 : OAI21_X1 port map( B1 => n629_port, B2 => n11355, A => n11120, ZN 
                           => N3676);
   U17269 : OAI21_X1 port map( B1 => n628_port, B2 => n11355, A => n11124, ZN 
                           => N3677);
   U17270 : OAI21_X1 port map( B1 => n627_port, B2 => n11355, A => n11128, ZN 
                           => N3678);
   U17271 : OAI21_X1 port map( B1 => n626_port, B2 => n11355, A => n11132, ZN 
                           => N3679);
   U17272 : OAI21_X1 port map( B1 => n625_port, B2 => n11354, A => n11136, ZN 
                           => N3680);
   U17273 : OAI21_X1 port map( B1 => n624_port, B2 => n11354, A => n11140, ZN 
                           => N3681);
   U17274 : OAI21_X1 port map( B1 => n623_port, B2 => n11354, A => n11144, ZN 
                           => N3682);
   U17275 : OAI21_X1 port map( B1 => n622_port, B2 => n11354, A => n11148, ZN 
                           => N3683);
   U17276 : OAI21_X1 port map( B1 => n621_port, B2 => n11354, A => n11152, ZN 
                           => N3684);
   U17277 : OAI21_X1 port map( B1 => n620_port, B2 => n11354, A => n11156, ZN 
                           => N3685);
   U17278 : OAI21_X1 port map( B1 => n619_port, B2 => n11354, A => n11160, ZN 
                           => N3686);
   U17279 : OAI21_X1 port map( B1 => n618_port, B2 => n11354, A => n11164, ZN 
                           => N3687);
   U17280 : OAI21_X1 port map( B1 => n617_port, B2 => n11354, A => n11168, ZN 
                           => N3688);
   U17281 : OAI21_X1 port map( B1 => n616_port, B2 => n11354, A => n11172, ZN 
                           => N3689);
   U17282 : OAI21_X1 port map( B1 => n615_port, B2 => n11354, A => n11176, ZN 
                           => N3690);
   U17283 : OAI21_X1 port map( B1 => n614_port, B2 => n11354, A => n11180, ZN 
                           => N3691);
   U17284 : OAI21_X1 port map( B1 => n613_port, B2 => n11353, A => n11184, ZN 
                           => N3692);
   U17285 : OAI21_X1 port map( B1 => n612_port, B2 => n11353, A => n11188, ZN 
                           => N3693);
   U17286 : OAI21_X1 port map( B1 => n611_port, B2 => n11353, A => n11192, ZN 
                           => N3694);
   U17287 : OAI21_X1 port map( B1 => n610_port, B2 => n11353, A => n11196, ZN 
                           => N3695);
   U17288 : OAI21_X1 port map( B1 => n609_port, B2 => n11353, A => n11200, ZN 
                           => N3696);
   U17289 : OAI21_X1 port map( B1 => n608_port, B2 => n11353, A => n11204, ZN 
                           => N3697);
   U17290 : OAI21_X1 port map( B1 => n607_port, B2 => n11353, A => n11208, ZN 
                           => N3698);
   U17291 : OAI21_X1 port map( B1 => n606_port, B2 => n11353, A => n11212, ZN 
                           => N3699);
   U17292 : OAI21_X1 port map( B1 => n605_port, B2 => n11353, A => n11216, ZN 
                           => N3700);
   U17293 : OAI21_X1 port map( B1 => n604_port, B2 => n11353, A => n11220, ZN 
                           => N3701);
   U17294 : OAI21_X1 port map( B1 => n603_port, B2 => n11353, A => n11224, ZN 
                           => N3702);
   U17295 : OAI21_X1 port map( B1 => n602_port, B2 => n11353, A => n11228, ZN 
                           => N3703);
   U17296 : OAI21_X1 port map( B1 => n601_port, B2 => n11352, A => n11232, ZN 
                           => N3704);
   U17297 : OAI21_X1 port map( B1 => n600_port, B2 => n11352, A => n11236, ZN 
                           => N3705);
   U17298 : OAI21_X1 port map( B1 => n599_port, B2 => n11352, A => n11240, ZN 
                           => N3706);
   U17299 : OAI21_X1 port map( B1 => n598_port, B2 => n11352, A => n11244, ZN 
                           => N3707);
   U17300 : OAI21_X1 port map( B1 => n597_port, B2 => n11352, A => n11248, ZN 
                           => N3708);
   U17301 : OAI21_X1 port map( B1 => n596_port, B2 => n11352, A => n11252, ZN 
                           => N3709);
   U17302 : OAI21_X1 port map( B1 => n595_port, B2 => n11352, A => n11256, ZN 
                           => N3710);
   U17303 : OAI21_X1 port map( B1 => n594_port, B2 => n11352, A => n11260, ZN 
                           => N3711);
   U17304 : OAI21_X1 port map( B1 => n593_port, B2 => n11352, A => n11264, ZN 
                           => N3712);
   U17305 : OAI21_X1 port map( B1 => n592_port, B2 => n11352, A => n11268, ZN 
                           => N3713);
   U17306 : OAI21_X1 port map( B1 => n591_port, B2 => n11352, A => n11272, ZN 
                           => N3714);
   U17307 : OAI21_X1 port map( B1 => n590_port, B2 => n11352, A => n11276, ZN 
                           => N3715);
   U17308 : OAI21_X1 port map( B1 => n589_port, B2 => n11351, A => n11280, ZN 
                           => N3716);
   U17309 : OAI21_X1 port map( B1 => n588_port, B2 => n11351, A => n11284, ZN 
                           => N3717);
   U17310 : OAI21_X1 port map( B1 => n587_port, B2 => n11351, A => n11288, ZN 
                           => N3718);
   U17311 : OAI21_X1 port map( B1 => n586_port, B2 => n11351, A => n11292, ZN 
                           => N3719);
   U17312 : OAI21_X1 port map( B1 => n585_port, B2 => n11351, A => n11296, ZN 
                           => N3720);
   U17313 : OAI21_X1 port map( B1 => n584_port, B2 => n11351, A => n11300, ZN 
                           => N3721);
   U17314 : OAI21_X1 port map( B1 => n583_port, B2 => n11351, A => n11304, ZN 
                           => N3722);
   U17315 : OAI21_X1 port map( B1 => n582_port, B2 => n11351, A => n11308, ZN 
                           => N3723);
   U17316 : OAI21_X1 port map( B1 => n581_port, B2 => n11351, A => n11312, ZN 
                           => N3724);
   U17317 : OAI21_X1 port map( B1 => n580_port, B2 => n11351, A => n11316, ZN 
                           => N3725);
   U17318 : OAI21_X1 port map( B1 => n579_port, B2 => n11351, A => n11320, ZN 
                           => N3726);
   U17319 : OAI21_X1 port map( B1 => n578_port, B2 => n11350, A => n11324, ZN 
                           => N3727);
   U17320 : OAI21_X1 port map( B1 => n577_port, B2 => n11350, A => n11328, ZN 
                           => N3728);
   U17321 : OAI21_X1 port map( B1 => n576_port, B2 => n11350, A => n11076, ZN 
                           => N3730);
   U17322 : OAI21_X1 port map( B1 => n575_port, B2 => n11350, A => n11080, ZN 
                           => N3731);
   U17323 : OAI21_X1 port map( B1 => n574_port, B2 => n11350, A => n11084, ZN 
                           => N3732);
   U17324 : OAI21_X1 port map( B1 => n573_port, B2 => n11350, A => n11088, ZN 
                           => N3733);
   U17325 : OAI21_X1 port map( B1 => n572_port, B2 => n11350, A => n11092, ZN 
                           => N3734);
   U17326 : OAI21_X1 port map( B1 => n571_port, B2 => n11350, A => n11096, ZN 
                           => N3735);
   U17327 : OAI21_X1 port map( B1 => n570_port, B2 => n11350, A => n11100, ZN 
                           => N3736);
   U17328 : OAI21_X1 port map( B1 => n569_port, B2 => n11350, A => n11104, ZN 
                           => N3737);
   U17329 : OAI21_X1 port map( B1 => n568_port, B2 => n11350, A => n11108, ZN 
                           => N3738);
   U17330 : OAI21_X1 port map( B1 => n567_port, B2 => n11350, A => n11112, ZN 
                           => N3739);
   U17331 : OAI21_X1 port map( B1 => n566_port, B2 => n11349, A => n11116, ZN 
                           => N3740);
   U17332 : OAI21_X1 port map( B1 => n565_port, B2 => n11349, A => n11120, ZN 
                           => N3741);
   U17333 : OAI21_X1 port map( B1 => n564_port, B2 => n11349, A => n11124, ZN 
                           => N3742);
   U17334 : OAI21_X1 port map( B1 => n563_port, B2 => n11349, A => n11128, ZN 
                           => N3743);
   U17335 : OAI21_X1 port map( B1 => n562_port, B2 => n11349, A => n11132, ZN 
                           => N3744);
   U17336 : OAI21_X1 port map( B1 => n561_port, B2 => n11349, A => n11136, ZN 
                           => N3745);
   U17337 : OAI21_X1 port map( B1 => n560_port, B2 => n11349, A => n11140, ZN 
                           => N3746);
   U17338 : OAI21_X1 port map( B1 => n559_port, B2 => n11349, A => n11144, ZN 
                           => N3747);
   U17339 : OAI21_X1 port map( B1 => n558_port, B2 => n11349, A => n11148, ZN 
                           => N3748);
   U17340 : OAI21_X1 port map( B1 => n557_port, B2 => n11349, A => n11152, ZN 
                           => N3749);
   U17341 : OAI21_X1 port map( B1 => n556_port, B2 => n11349, A => n11156, ZN 
                           => N3750);
   U17342 : OAI21_X1 port map( B1 => n555_port, B2 => n11349, A => n11160, ZN 
                           => N3751);
   U17343 : OAI21_X1 port map( B1 => n554_port, B2 => n11348, A => n11164, ZN 
                           => N3752);
   U17344 : OAI21_X1 port map( B1 => n553_port, B2 => n11348, A => n11168, ZN 
                           => N3753);
   U17345 : OAI21_X1 port map( B1 => n552_port, B2 => n11348, A => n11172, ZN 
                           => N3754);
   U17346 : OAI21_X1 port map( B1 => n551_port, B2 => n11348, A => n11176, ZN 
                           => N3755);
   U17347 : OAI21_X1 port map( B1 => n550_port, B2 => n11348, A => n11180, ZN 
                           => N3756);
   U17348 : OAI21_X1 port map( B1 => n549_port, B2 => n11348, A => n11184, ZN 
                           => N3757);
   U17349 : OAI21_X1 port map( B1 => n548_port, B2 => n11348, A => n11188, ZN 
                           => N3758);
   U17350 : OAI21_X1 port map( B1 => n547_port, B2 => n11348, A => n11192, ZN 
                           => N3759);
   U17351 : OAI21_X1 port map( B1 => n546_port, B2 => n11348, A => n11196, ZN 
                           => N3760);
   U17352 : OAI21_X1 port map( B1 => n545_port, B2 => n11348, A => n11200, ZN 
                           => N3761);
   U17353 : OAI21_X1 port map( B1 => n544_port, B2 => n11348, A => n11204, ZN 
                           => N3762);
   U17354 : OAI21_X1 port map( B1 => n543_port, B2 => n11348, A => n11208, ZN 
                           => N3763);
   U17355 : OAI21_X1 port map( B1 => n542_port, B2 => n11347, A => n11212, ZN 
                           => N3764);
   U17356 : OAI21_X1 port map( B1 => n541_port, B2 => n11347, A => n11216, ZN 
                           => N3765);
   U17357 : OAI21_X1 port map( B1 => n540_port, B2 => n11347, A => n11220, ZN 
                           => N3766);
   U17358 : OAI21_X1 port map( B1 => n539_port, B2 => n11347, A => n11224, ZN 
                           => N3767);
   U17359 : OAI21_X1 port map( B1 => n538_port, B2 => n11347, A => n11228, ZN 
                           => N3768);
   U17360 : OAI21_X1 port map( B1 => n537_port, B2 => n11347, A => n11232, ZN 
                           => N3769);
   U17361 : OAI21_X1 port map( B1 => n536_port, B2 => n11347, A => n11236, ZN 
                           => N3770);
   U17362 : OAI21_X1 port map( B1 => n535_port, B2 => n11347, A => n11240, ZN 
                           => N3771);
   U17363 : OAI21_X1 port map( B1 => n534_port, B2 => n11347, A => n11244, ZN 
                           => N3772);
   U17364 : OAI21_X1 port map( B1 => n533_port, B2 => n11347, A => n11248, ZN 
                           => N3773);
   U17365 : OAI21_X1 port map( B1 => n532_port, B2 => n11347, A => n11252, ZN 
                           => N3774);
   U17366 : OAI21_X1 port map( B1 => n531_port, B2 => n11347, A => n11256, ZN 
                           => N3775);
   U17367 : OAI21_X1 port map( B1 => n530_port, B2 => n11346, A => n11260, ZN 
                           => N3776);
   U17368 : OAI21_X1 port map( B1 => n529_port, B2 => n11346, A => n11264, ZN 
                           => N3777);
   U17369 : OAI21_X1 port map( B1 => n528_port, B2 => n11346, A => n11268, ZN 
                           => N3778);
   U17370 : OAI21_X1 port map( B1 => n527_port, B2 => n11346, A => n11272, ZN 
                           => N3779);
   U17371 : OAI21_X1 port map( B1 => n526_port, B2 => n11346, A => n11276, ZN 
                           => N3780);
   U17372 : OAI21_X1 port map( B1 => n525_port, B2 => n11346, A => n11280, ZN 
                           => N3781);
   U17373 : OAI21_X1 port map( B1 => n524_port, B2 => n11346, A => n11284, ZN 
                           => N3782);
   U17374 : OAI21_X1 port map( B1 => n523_port, B2 => n11346, A => n11288, ZN 
                           => N3783);
   U17375 : OAI21_X1 port map( B1 => n522_port, B2 => n11346, A => n11292, ZN 
                           => N3784);
   U17376 : OAI21_X1 port map( B1 => n521_port, B2 => n11346, A => n11296, ZN 
                           => N3785);
   U17377 : OAI21_X1 port map( B1 => n520_port, B2 => n11346, A => n11300, ZN 
                           => N3786);
   U17378 : OAI21_X1 port map( B1 => n519_port, B2 => n11351, A => n11304, ZN 
                           => N3787);
   U17379 : OAI21_X1 port map( B1 => n518_port, B2 => n11356, A => n11308, ZN 
                           => N3788);
   U17380 : OAI21_X1 port map( B1 => n517_port, B2 => n11410, A => n11312, ZN 
                           => N3789);
   U17381 : OAI21_X1 port map( B1 => n516_port, B2 => n11410, A => n11316, ZN 
                           => N3790);
   U17382 : OAI21_X1 port map( B1 => n515_port, B2 => n11410, A => n11320, ZN 
                           => N3791);
   U17383 : OAI21_X1 port map( B1 => n514_port, B2 => n11410, A => n11324, ZN 
                           => N3792);
   U17384 : OAI21_X1 port map( B1 => n513_port, B2 => n11410, A => n11328, ZN 
                           => N3793);
   U17385 : OAI21_X1 port map( B1 => n512_port, B2 => n11410, A => n11077, ZN 
                           => N3795);
   U17386 : OAI21_X1 port map( B1 => n511_port, B2 => n11410, A => n11081, ZN 
                           => N3796);
   U17387 : OAI21_X1 port map( B1 => n510_port, B2 => n11409, A => n11085, ZN 
                           => N3797);
   U17388 : OAI21_X1 port map( B1 => n509_port, B2 => n11409, A => n11089, ZN 
                           => N3798);
   U17389 : OAI21_X1 port map( B1 => n508_port, B2 => n11409, A => n11093, ZN 
                           => N3799);
   U17390 : OAI21_X1 port map( B1 => n507_port, B2 => n11409, A => n11097, ZN 
                           => N3800);
   U17391 : OAI21_X1 port map( B1 => n506_port, B2 => n11409, A => n11101, ZN 
                           => N3801);
   U17392 : OAI21_X1 port map( B1 => n505_port, B2 => n11409, A => n11105, ZN 
                           => N3802);
   U17393 : OAI21_X1 port map( B1 => n504_port, B2 => n11409, A => n11109, ZN 
                           => N3803);
   U17394 : OAI21_X1 port map( B1 => n503_port, B2 => n11409, A => n11113, ZN 
                           => N3804);
   U17395 : OAI21_X1 port map( B1 => n502_port, B2 => n11409, A => n11117, ZN 
                           => N3805);
   U17396 : OAI21_X1 port map( B1 => n501_port, B2 => n11409, A => n11121, ZN 
                           => N3806);
   U17397 : OAI21_X1 port map( B1 => n500_port, B2 => n11409, A => n11125, ZN 
                           => N3807);
   U17398 : OAI21_X1 port map( B1 => n499_port, B2 => n11409, A => n11129, ZN 
                           => N3808);
   U17399 : OAI21_X1 port map( B1 => n498_port, B2 => n11408, A => n11133, ZN 
                           => N3809);
   U17400 : OAI21_X1 port map( B1 => n497_port, B2 => n11408, A => n11137, ZN 
                           => N3810);
   U17401 : OAI21_X1 port map( B1 => n496_port, B2 => n11408, A => n11141, ZN 
                           => N3811);
   U17402 : OAI21_X1 port map( B1 => n495_port, B2 => n11408, A => n11145, ZN 
                           => N3812);
   U17403 : OAI21_X1 port map( B1 => n494_port, B2 => n11408, A => n11149, ZN 
                           => N3813);
   U17404 : OAI21_X1 port map( B1 => n493_port, B2 => n11408, A => n11153, ZN 
                           => N3814);
   U17405 : OAI21_X1 port map( B1 => n492_port, B2 => n11408, A => n11157, ZN 
                           => N3815);
   U17406 : OAI21_X1 port map( B1 => n491_port, B2 => n11408, A => n11161, ZN 
                           => N3816);
   U17407 : OAI21_X1 port map( B1 => n490_port, B2 => n11408, A => n11165, ZN 
                           => N3817);
   U17408 : OAI21_X1 port map( B1 => n489_port, B2 => n11408, A => n11169, ZN 
                           => N3818);
   U17409 : OAI21_X1 port map( B1 => n488_port, B2 => n11408, A => n11173, ZN 
                           => N3819);
   U17410 : OAI21_X1 port map( B1 => n487_port, B2 => n11408, A => n11177, ZN 
                           => N3820);
   U17411 : OAI21_X1 port map( B1 => n486_port, B2 => n11407, A => n11181, ZN 
                           => N3821);
   U17412 : OAI21_X1 port map( B1 => n485_port, B2 => n11407, A => n11185, ZN 
                           => N3822);
   U17413 : OAI21_X1 port map( B1 => n484_port, B2 => n11407, A => n11189, ZN 
                           => N3823);
   U17414 : OAI21_X1 port map( B1 => n483_port, B2 => n11407, A => n11193, ZN 
                           => N3824);
   U17415 : OAI21_X1 port map( B1 => n482_port, B2 => n11407, A => n11197, ZN 
                           => N3825);
   U17416 : OAI21_X1 port map( B1 => n481_port, B2 => n11407, A => n11201, ZN 
                           => N3826);
   U17417 : OAI21_X1 port map( B1 => n480_port, B2 => n11407, A => n11205, ZN 
                           => N3827);
   U17418 : OAI21_X1 port map( B1 => n479_port, B2 => n11407, A => n11209, ZN 
                           => N3828);
   U17419 : OAI21_X1 port map( B1 => n478_port, B2 => n11407, A => n11213, ZN 
                           => N3829);
   U17420 : OAI21_X1 port map( B1 => n477_port, B2 => n11407, A => n11217, ZN 
                           => N3830);
   U17421 : OAI21_X1 port map( B1 => n476_port, B2 => n11407, A => n11221, ZN 
                           => N3831);
   U17422 : OAI21_X1 port map( B1 => n475_port, B2 => n11407, A => n11225, ZN 
                           => N3832);
   U17423 : OAI21_X1 port map( B1 => n474_port, B2 => n11406, A => n11229, ZN 
                           => N3833);
   U17424 : OAI21_X1 port map( B1 => n473_port, B2 => n11406, A => n11233, ZN 
                           => N3834);
   U17425 : OAI21_X1 port map( B1 => n472_port, B2 => n11406, A => n11237, ZN 
                           => N3835);
   U17426 : OAI21_X1 port map( B1 => n471_port, B2 => n11406, A => n11241, ZN 
                           => N3836);
   U17427 : OAI21_X1 port map( B1 => n470_port, B2 => n11406, A => n11245, ZN 
                           => N3837);
   U17428 : OAI21_X1 port map( B1 => n469_port, B2 => n11406, A => n11249, ZN 
                           => N3838);
   U17429 : OAI21_X1 port map( B1 => n468_port, B2 => n11406, A => n11253, ZN 
                           => N3839);
   U17430 : OAI21_X1 port map( B1 => n467_port, B2 => n11406, A => n11257, ZN 
                           => N3840);
   U17431 : OAI21_X1 port map( B1 => n466_port, B2 => n11406, A => n11261, ZN 
                           => N3841);
   U17432 : OAI21_X1 port map( B1 => n465_port, B2 => n11406, A => n11265, ZN 
                           => N3842);
   U17433 : OAI21_X1 port map( B1 => n464_port, B2 => n11406, A => n11269, ZN 
                           => N3843);
   U17434 : OAI21_X1 port map( B1 => n463_port, B2 => n11406, A => n11273, ZN 
                           => N3844);
   U17435 : OAI21_X1 port map( B1 => n462_port, B2 => n11405, A => n11277, ZN 
                           => N3845);
   U17436 : OAI21_X1 port map( B1 => n461_port, B2 => n11405, A => n11281, ZN 
                           => N3846);
   U17437 : OAI21_X1 port map( B1 => n460_port, B2 => n11405, A => n11285, ZN 
                           => N3847);
   U17438 : OAI21_X1 port map( B1 => n459_port, B2 => n11405, A => n11289, ZN 
                           => N3848);
   U17439 : OAI21_X1 port map( B1 => n458_port, B2 => n11405, A => n11293, ZN 
                           => N3849);
   U17440 : OAI21_X1 port map( B1 => n457_port, B2 => n11405, A => n11297, ZN 
                           => N3850);
   U17441 : OAI21_X1 port map( B1 => n456_port, B2 => n11405, A => n11301, ZN 
                           => N3851);
   U17442 : OAI21_X1 port map( B1 => n455_port, B2 => n11405, A => n11305, ZN 
                           => N3852);
   U17443 : OAI21_X1 port map( B1 => n454_port, B2 => n11405, A => n11309, ZN 
                           => N3853);
   U17444 : OAI21_X1 port map( B1 => n453_port, B2 => n11405, A => n11313, ZN 
                           => N3854);
   U17445 : OAI21_X1 port map( B1 => n452_port, B2 => n11405, A => n11317, ZN 
                           => N3855);
   U17446 : OAI21_X1 port map( B1 => n451_port, B2 => n11404, A => n11321, ZN 
                           => N3856);
   U17447 : OAI21_X1 port map( B1 => n450_port, B2 => n11404, A => n11325, ZN 
                           => N3857);
   U17448 : OAI21_X1 port map( B1 => n449_port, B2 => n11404, A => n11329, ZN 
                           => N3858);
   U17449 : OAI21_X1 port map( B1 => n448_port, B2 => n11404, A => n11077, ZN 
                           => N3860);
   U17450 : OAI21_X1 port map( B1 => n447_port, B2 => n11404, A => n11081, ZN 
                           => N3861);
   U17451 : OAI21_X1 port map( B1 => n446_port, B2 => n11404, A => n11085, ZN 
                           => N3862);
   U17452 : OAI21_X1 port map( B1 => n445_port, B2 => n11404, A => n11089, ZN 
                           => N3863);
   U17453 : OAI21_X1 port map( B1 => n444_port, B2 => n11404, A => n11093, ZN 
                           => N3864);
   U17454 : OAI21_X1 port map( B1 => n443_port, B2 => n11404, A => n11097, ZN 
                           => N3865);
   U17455 : OAI21_X1 port map( B1 => n442_port, B2 => n11404, A => n11101, ZN 
                           => N3866);
   U17456 : OAI21_X1 port map( B1 => n441_port, B2 => n11404, A => n11105, ZN 
                           => N3867);
   U17457 : OAI21_X1 port map( B1 => n440_port, B2 => n11404, A => n11109, ZN 
                           => N3868);
   U17458 : OAI21_X1 port map( B1 => n439_port, B2 => n11403, A => n11113, ZN 
                           => N3869);
   U17459 : OAI21_X1 port map( B1 => n438_port, B2 => n11403, A => n11117, ZN 
                           => N3870);
   U17460 : OAI21_X1 port map( B1 => n437_port, B2 => n11403, A => n11121, ZN 
                           => N3871);
   U17461 : OAI21_X1 port map( B1 => n436_port, B2 => n11403, A => n11125, ZN 
                           => N3872);
   U17462 : OAI21_X1 port map( B1 => n435_port, B2 => n11403, A => n11129, ZN 
                           => N3873);
   U17463 : OAI21_X1 port map( B1 => n434_port, B2 => n11403, A => n11133, ZN 
                           => N3874);
   U17464 : OAI21_X1 port map( B1 => n433_port, B2 => n11403, A => n11137, ZN 
                           => N3875);
   U17465 : OAI21_X1 port map( B1 => n432_port, B2 => n11403, A => n11141, ZN 
                           => N3876);
   U17466 : OAI21_X1 port map( B1 => n431_port, B2 => n11403, A => n11145, ZN 
                           => N3877);
   U17467 : OAI21_X1 port map( B1 => n430_port, B2 => n11403, A => n11149, ZN 
                           => N3878);
   U17468 : OAI21_X1 port map( B1 => n429_port, B2 => n11403, A => n11153, ZN 
                           => N3879);
   U17469 : OAI21_X1 port map( B1 => n428_port, B2 => n11403, A => n11157, ZN 
                           => N3880);
   U17470 : OAI21_X1 port map( B1 => n427_port, B2 => n11402, A => n11161, ZN 
                           => N3881);
   U17471 : OAI21_X1 port map( B1 => n426_port, B2 => n11402, A => n11165, ZN 
                           => N3882);
   U17472 : OAI21_X1 port map( B1 => n425_port, B2 => n11402, A => n11169, ZN 
                           => N3883);
   U17473 : OAI21_X1 port map( B1 => n424_port, B2 => n11402, A => n11173, ZN 
                           => N3884);
   U17474 : OAI21_X1 port map( B1 => n423_port, B2 => n11402, A => n11177, ZN 
                           => N3885);
   U17475 : OAI21_X1 port map( B1 => n422_port, B2 => n11402, A => n11181, ZN 
                           => N3886);
   U17476 : OAI21_X1 port map( B1 => n421_port, B2 => n11402, A => n11185, ZN 
                           => N3887);
   U17477 : OAI21_X1 port map( B1 => n420_port, B2 => n11402, A => n11189, ZN 
                           => N3888);
   U17478 : OAI21_X1 port map( B1 => n419_port, B2 => n11402, A => n11193, ZN 
                           => N3889);
   U17479 : OAI21_X1 port map( B1 => n418_port, B2 => n11402, A => n11197, ZN 
                           => N3890);
   U17480 : OAI21_X1 port map( B1 => n417_port, B2 => n11402, A => n11201, ZN 
                           => N3891);
   U17481 : OAI21_X1 port map( B1 => n416_port, B2 => n11402, A => n11205, ZN 
                           => N3892);
   U17482 : OAI21_X1 port map( B1 => n415_port, B2 => n11401, A => n11209, ZN 
                           => N3893);
   U17483 : OAI21_X1 port map( B1 => n414_port, B2 => n11401, A => n11213, ZN 
                           => N3894);
   U17484 : OAI21_X1 port map( B1 => n413_port, B2 => n11401, A => n11217, ZN 
                           => N3895);
   U17485 : OAI21_X1 port map( B1 => n412_port, B2 => n11401, A => n11221, ZN 
                           => N3896);
   U17486 : OAI21_X1 port map( B1 => n411_port, B2 => n11401, A => n11225, ZN 
                           => N3897);
   U17487 : OAI21_X1 port map( B1 => n410_port, B2 => n11401, A => n11229, ZN 
                           => N3898);
   U17488 : OAI21_X1 port map( B1 => n409_port, B2 => n11401, A => n11233, ZN 
                           => N3899);
   U17489 : OAI21_X1 port map( B1 => n408_port, B2 => n11401, A => n11237, ZN 
                           => N3900);
   U17490 : OAI21_X1 port map( B1 => n407_port, B2 => n11401, A => n11241, ZN 
                           => N3901);
   U17491 : OAI21_X1 port map( B1 => n406_port, B2 => n11401, A => n11245, ZN 
                           => N3902);
   U17492 : OAI21_X1 port map( B1 => n405_port, B2 => n11401, A => n11249, ZN 
                           => N3903);
   U17493 : OAI21_X1 port map( B1 => n404_port, B2 => n11401, A => n11253, ZN 
                           => N3904);
   U17494 : OAI21_X1 port map( B1 => n403_port, B2 => n11400, A => n11257, ZN 
                           => N3905);
   U17495 : OAI21_X1 port map( B1 => n402_port, B2 => n11400, A => n11261, ZN 
                           => N3906);
   U17496 : OAI21_X1 port map( B1 => n401_port, B2 => n11400, A => n11265, ZN 
                           => N3907);
   U17497 : OAI21_X1 port map( B1 => n400_port, B2 => n11400, A => n11269, ZN 
                           => N3908);
   U17498 : OAI21_X1 port map( B1 => n399_port, B2 => n11400, A => n11273, ZN 
                           => N3909);
   U17499 : OAI21_X1 port map( B1 => n398_port, B2 => n11400, A => n11277, ZN 
                           => N3910);
   U17500 : OAI21_X1 port map( B1 => n397_port, B2 => n11400, A => n11281, ZN 
                           => N3911);
   U17501 : OAI21_X1 port map( B1 => n396_port, B2 => n11400, A => n11285, ZN 
                           => N3912);
   U17502 : OAI21_X1 port map( B1 => n395_port, B2 => n11400, A => n11289, ZN 
                           => N3913);
   U17503 : OAI21_X1 port map( B1 => n394_port, B2 => n11400, A => n11293, ZN 
                           => N3914);
   U17504 : OAI21_X1 port map( B1 => n393_port, B2 => n11400, A => n11297, ZN 
                           => N3915);
   U17505 : OAI21_X1 port map( B1 => n392_port, B2 => n11400, A => n11301, ZN 
                           => N3916);
   U17506 : OAI21_X1 port map( B1 => n391_port, B2 => n11399, A => n11305, ZN 
                           => N3917);
   U17507 : OAI21_X1 port map( B1 => n390_port, B2 => n11399, A => n11309, ZN 
                           => N3918);
   U17508 : OAI21_X1 port map( B1 => n389_port, B2 => n11405, A => n11313, ZN 
                           => N3919);
   U17509 : OAI21_X1 port map( B1 => n388_port, B2 => n11421, A => n11317, ZN 
                           => N3920);
   U17510 : OAI21_X1 port map( B1 => n387_port, B2 => n11421, A => n11321, ZN 
                           => N3921);
   U17511 : OAI21_X1 port map( B1 => n386_port, B2 => n11421, A => n11325, ZN 
                           => N3922);
   U17512 : OAI21_X1 port map( B1 => n385_port, B2 => n11420, A => n11329, ZN 
                           => N3923);
   U17513 : OAI21_X1 port map( B1 => n384_port, B2 => n11420, A => n11077, ZN 
                           => N3925);
   U17514 : OAI21_X1 port map( B1 => n383_port, B2 => n11420, A => n11081, ZN 
                           => N3926);
   U17515 : OAI21_X1 port map( B1 => n382_port, B2 => n11420, A => n11085, ZN 
                           => N3927);
   U17516 : OAI21_X1 port map( B1 => n381_port, B2 => n11420, A => n11089, ZN 
                           => N3928);
   U17517 : OAI21_X1 port map( B1 => n380_port, B2 => n11420, A => n11093, ZN 
                           => N3929);
   U17518 : OAI21_X1 port map( B1 => n379_port, B2 => n11420, A => n11097, ZN 
                           => N3930);
   U17519 : OAI21_X1 port map( B1 => n378_port, B2 => n11420, A => n11101, ZN 
                           => N3931);
   U17520 : OAI21_X1 port map( B1 => n377_port, B2 => n11420, A => n11105, ZN 
                           => N3932);
   U17521 : OAI21_X1 port map( B1 => n376_port, B2 => n11420, A => n11109, ZN 
                           => N3933);
   U17522 : OAI21_X1 port map( B1 => n375_port, B2 => n11420, A => n11113, ZN 
                           => N3934);
   U17523 : OAI21_X1 port map( B1 => n374_port, B2 => n11420, A => n11117, ZN 
                           => N3935);
   U17524 : OAI21_X1 port map( B1 => n373_port, B2 => n11419, A => n11121, ZN 
                           => N3936);
   U17525 : OAI21_X1 port map( B1 => n372_port, B2 => n11419, A => n11125, ZN 
                           => N3937);
   U17526 : OAI21_X1 port map( B1 => n371_port, B2 => n11419, A => n11129, ZN 
                           => N3938);
   U17527 : OAI21_X1 port map( B1 => n370_port, B2 => n11419, A => n11133, ZN 
                           => N3939);
   U17528 : OAI21_X1 port map( B1 => n369_port, B2 => n11419, A => n11137, ZN 
                           => N3940);
   U17529 : OAI21_X1 port map( B1 => n368_port, B2 => n11419, A => n11141, ZN 
                           => N3941);
   U17530 : OAI21_X1 port map( B1 => n367_port, B2 => n11419, A => n11145, ZN 
                           => N3942);
   U17531 : OAI21_X1 port map( B1 => n366_port, B2 => n11419, A => n11149, ZN 
                           => N3943);
   U17532 : OAI21_X1 port map( B1 => n365_port, B2 => n11419, A => n11153, ZN 
                           => N3944);
   U17533 : OAI21_X1 port map( B1 => n364_port, B2 => n11419, A => n11157, ZN 
                           => N3945);
   U17534 : OAI21_X1 port map( B1 => n363_port, B2 => n11419, A => n11161, ZN 
                           => N3946);
   U17535 : OAI21_X1 port map( B1 => n362_port, B2 => n11419, A => n11165, ZN 
                           => N3947);
   U17536 : OAI21_X1 port map( B1 => n361_port, B2 => n11418, A => n11169, ZN 
                           => N3948);
   U17537 : OAI21_X1 port map( B1 => n360_port, B2 => n11418, A => n11173, ZN 
                           => N3949);
   U17538 : OAI21_X1 port map( B1 => n359_port, B2 => n11418, A => n11177, ZN 
                           => N3950);
   U17539 : OAI21_X1 port map( B1 => n358_port, B2 => n11418, A => n11181, ZN 
                           => N3951);
   U17540 : OAI21_X1 port map( B1 => n357_port, B2 => n11418, A => n11185, ZN 
                           => N3952);
   U17541 : OAI21_X1 port map( B1 => n356_port, B2 => n11418, A => n11189, ZN 
                           => N3953);
   U17542 : OAI21_X1 port map( B1 => n355_port, B2 => n11418, A => n11193, ZN 
                           => N3954);
   U17543 : OAI21_X1 port map( B1 => n354_port, B2 => n11418, A => n11197, ZN 
                           => N3955);
   U17544 : OAI21_X1 port map( B1 => n353_port, B2 => n11418, A => n11201, ZN 
                           => N3956);
   U17545 : OAI21_X1 port map( B1 => n352_port, B2 => n11418, A => n11205, ZN 
                           => N3957);
   U17546 : OAI21_X1 port map( B1 => n351_port, B2 => n11418, A => n11209, ZN 
                           => N3958);
   U17547 : OAI21_X1 port map( B1 => n350_port, B2 => n11418, A => n11213, ZN 
                           => N3959);
   U17548 : OAI21_X1 port map( B1 => n349_port, B2 => n11417, A => n11217, ZN 
                           => N3960);
   U17549 : OAI21_X1 port map( B1 => n348_port, B2 => n11417, A => n11221, ZN 
                           => N3961);
   U17550 : OAI21_X1 port map( B1 => n347_port, B2 => n11417, A => n11225, ZN 
                           => N3962);
   U17551 : OAI21_X1 port map( B1 => n346_port, B2 => n11417, A => n11229, ZN 
                           => N3963);
   U17552 : OAI21_X1 port map( B1 => n345_port, B2 => n11417, A => n11233, ZN 
                           => N3964);
   U17553 : OAI21_X1 port map( B1 => n344_port, B2 => n11417, A => n11237, ZN 
                           => N3965);
   U17554 : OAI21_X1 port map( B1 => n343_port, B2 => n11417, A => n11241, ZN 
                           => N3966);
   U17555 : OAI21_X1 port map( B1 => n342_port, B2 => n11417, A => n11245, ZN 
                           => N3967);
   U17556 : OAI21_X1 port map( B1 => n341_port, B2 => n11417, A => n11249, ZN 
                           => N3968);
   U17557 : OAI21_X1 port map( B1 => n340_port, B2 => n11417, A => n11253, ZN 
                           => N3969);
   U17558 : OAI21_X1 port map( B1 => n339_port, B2 => n11417, A => n11257, ZN 
                           => N3970);
   U17559 : OAI21_X1 port map( B1 => n338_port, B2 => n11417, A => n11261, ZN 
                           => N3971);
   U17560 : OAI21_X1 port map( B1 => n337_port, B2 => n11416, A => n11265, ZN 
                           => N3972);
   U17561 : OAI21_X1 port map( B1 => n336_port, B2 => n11416, A => n11269, ZN 
                           => N3973);
   U17562 : OAI21_X1 port map( B1 => n335_port, B2 => n11416, A => n11273, ZN 
                           => N3974);
   U17563 : OAI21_X1 port map( B1 => n334_port, B2 => n11416, A => n11277, ZN 
                           => N3975);
   U17564 : OAI21_X1 port map( B1 => n333_port, B2 => n11416, A => n11281, ZN 
                           => N3976);
   U17565 : OAI21_X1 port map( B1 => n332_port, B2 => n11416, A => n11285, ZN 
                           => N3977);
   U17566 : OAI21_X1 port map( B1 => n331_port, B2 => n11416, A => n11289, ZN 
                           => N3978);
   U17567 : OAI21_X1 port map( B1 => n330_port, B2 => n11416, A => n11293, ZN 
                           => N3979);
   U17568 : OAI21_X1 port map( B1 => n329_port, B2 => n11416, A => n11297, ZN 
                           => N3980);
   U17569 : OAI21_X1 port map( B1 => n328_port, B2 => n11416, A => n11301, ZN 
                           => N3981);
   U17570 : OAI21_X1 port map( B1 => n327_port, B2 => n11416, A => n11305, ZN 
                           => N3982);
   U17571 : OAI21_X1 port map( B1 => n326_port, B2 => n11416, A => n11309, ZN 
                           => N3983);
   U17572 : OAI21_X1 port map( B1 => n325_port, B2 => n11415, A => n11313, ZN 
                           => N3984);
   U17573 : OAI21_X1 port map( B1 => n324_port, B2 => n11415, A => n11317, ZN 
                           => N3985);
   U17574 : OAI21_X1 port map( B1 => n323_port, B2 => n11415, A => n11321, ZN 
                           => N3986);
   U17575 : OAI21_X1 port map( B1 => n322_port, B2 => n11415, A => n11325, ZN 
                           => N3987);
   U17576 : OAI21_X1 port map( B1 => n321_port, B2 => n11415, A => n11329, ZN 
                           => N3988);
   U17577 : OAI21_X1 port map( B1 => n320_port, B2 => n11415, A => n11077, ZN 
                           => N3990);
   U17578 : OAI21_X1 port map( B1 => n319_port, B2 => n11415, A => n11081, ZN 
                           => N3991);
   U17579 : OAI21_X1 port map( B1 => n318_port, B2 => n11415, A => n11085, ZN 
                           => N3992);
   U17580 : OAI21_X1 port map( B1 => n317_port, B2 => n11415, A => n11089, ZN 
                           => N3993);
   U17581 : OAI21_X1 port map( B1 => n316_port, B2 => n11415, A => n11093, ZN 
                           => N3994);
   U17582 : OAI21_X1 port map( B1 => n315_port, B2 => n11415, A => n11097, ZN 
                           => N3995);
   U17583 : OAI21_X1 port map( B1 => n314_port, B2 => n11414, A => n11101, ZN 
                           => N3996);
   U17584 : OAI21_X1 port map( B1 => n313_port, B2 => n11414, A => n11105, ZN 
                           => N3997);
   U17585 : OAI21_X1 port map( B1 => n312_port, B2 => n11414, A => n11109, ZN 
                           => N3998);
   U17586 : OAI21_X1 port map( B1 => n311_port, B2 => n11414, A => n11113, ZN 
                           => N3999);
   U17587 : OAI21_X1 port map( B1 => n310_port, B2 => n11414, A => n11117, ZN 
                           => N4000);
   U17588 : OAI21_X1 port map( B1 => n309_port, B2 => n11414, A => n11121, ZN 
                           => N4001);
   U17589 : OAI21_X1 port map( B1 => n308_port, B2 => n11414, A => n11125, ZN 
                           => N4002);
   U17590 : OAI21_X1 port map( B1 => n307_port, B2 => n11414, A => n11129, ZN 
                           => N4003);
   U17591 : OAI21_X1 port map( B1 => n306_port, B2 => n11414, A => n11133, ZN 
                           => N4004);
   U17592 : OAI21_X1 port map( B1 => n305_port, B2 => n11414, A => n11137, ZN 
                           => N4005);
   U17593 : OAI21_X1 port map( B1 => n304_port, B2 => n11414, A => n11141, ZN 
                           => N4006);
   U17594 : OAI21_X1 port map( B1 => n303_port, B2 => n11414, A => n11145, ZN 
                           => N4007);
   U17595 : OAI21_X1 port map( B1 => n302_port, B2 => n11413, A => n11149, ZN 
                           => N4008);
   U17596 : OAI21_X1 port map( B1 => n301_port, B2 => n11413, A => n11153, ZN 
                           => N4009);
   U17597 : OAI21_X1 port map( B1 => n300_port, B2 => n11413, A => n11157, ZN 
                           => N4010);
   U17598 : OAI21_X1 port map( B1 => n299_port, B2 => n11413, A => n11161, ZN 
                           => N4011);
   U17599 : OAI21_X1 port map( B1 => n298_port, B2 => n11413, A => n11165, ZN 
                           => N4012);
   U17600 : OAI21_X1 port map( B1 => n297_port, B2 => n11413, A => n11169, ZN 
                           => N4013);
   U17601 : OAI21_X1 port map( B1 => n296_port, B2 => n11413, A => n11173, ZN 
                           => N4014);
   U17602 : OAI21_X1 port map( B1 => n295_port, B2 => n11413, A => n11177, ZN 
                           => N4015);
   U17603 : OAI21_X1 port map( B1 => n294_port, B2 => n11413, A => n11181, ZN 
                           => N4016);
   U17604 : OAI21_X1 port map( B1 => n293_port, B2 => n11413, A => n11185, ZN 
                           => N4017);
   U17605 : OAI21_X1 port map( B1 => n292_port, B2 => n11413, A => n11189, ZN 
                           => N4018);
   U17606 : OAI21_X1 port map( B1 => n291_port, B2 => n11413, A => n11193, ZN 
                           => N4019);
   U17607 : OAI21_X1 port map( B1 => n290_port, B2 => n11412, A => n11197, ZN 
                           => N4020);
   U17608 : OAI21_X1 port map( B1 => n289_port, B2 => n11412, A => n11201, ZN 
                           => N4021);
   U17609 : OAI21_X1 port map( B1 => n288_port, B2 => n11412, A => n11205, ZN 
                           => N4022);
   U17610 : OAI21_X1 port map( B1 => n287_port, B2 => n11412, A => n11209, ZN 
                           => N4023);
   U17611 : OAI21_X1 port map( B1 => n286_port, B2 => n11412, A => n11213, ZN 
                           => N4024);
   U17612 : OAI21_X1 port map( B1 => n285_port, B2 => n11412, A => n11217, ZN 
                           => N4025);
   U17613 : OAI21_X1 port map( B1 => n284_port, B2 => n11412, A => n11221, ZN 
                           => N4026);
   U17614 : OAI21_X1 port map( B1 => n283_port, B2 => n11412, A => n11225, ZN 
                           => N4027);
   U17615 : OAI21_X1 port map( B1 => n282_port, B2 => n11412, A => n11229, ZN 
                           => N4028);
   U17616 : OAI21_X1 port map( B1 => n281_port, B2 => n11412, A => n11233, ZN 
                           => N4029);
   U17617 : OAI21_X1 port map( B1 => n280_port, B2 => n11412, A => n11237, ZN 
                           => N4030);
   U17618 : OAI21_X1 port map( B1 => n279_port, B2 => n11412, A => n11241, ZN 
                           => N4031);
   U17619 : OAI21_X1 port map( B1 => n278_port, B2 => n11411, A => n11245, ZN 
                           => N4032);
   U17620 : OAI21_X1 port map( B1 => n277_port, B2 => n11411, A => n11249, ZN 
                           => N4033);
   U17621 : OAI21_X1 port map( B1 => n276_port, B2 => n11411, A => n11253, ZN 
                           => N4034);
   U17622 : OAI21_X1 port map( B1 => n275_port, B2 => n11411, A => n11257, ZN 
                           => N4035);
   U17623 : OAI21_X1 port map( B1 => n274_port, B2 => n11411, A => n11261, ZN 
                           => N4036);
   U17624 : OAI21_X1 port map( B1 => n273_port, B2 => n11411, A => n11265, ZN 
                           => N4037);
   U17625 : OAI21_X1 port map( B1 => n272_port, B2 => n11411, A => n11269, ZN 
                           => N4038);
   U17626 : OAI21_X1 port map( B1 => n271_port, B2 => n11411, A => n11273, ZN 
                           => N4039);
   U17627 : OAI21_X1 port map( B1 => n270_port, B2 => n11411, A => n11277, ZN 
                           => N4040);
   U17628 : OAI21_X1 port map( B1 => n269_port, B2 => n11411, A => n11281, ZN 
                           => N4041);
   U17629 : OAI21_X1 port map( B1 => n268_port, B2 => n11411, A => n11285, ZN 
                           => N4042);
   U17630 : OAI21_X1 port map( B1 => n267_port, B2 => n11411, A => n11289, ZN 
                           => N4043);
   U17631 : OAI21_X1 port map( B1 => n266_port, B2 => n11410, A => n11293, ZN 
                           => N4044);
   U17632 : OAI21_X1 port map( B1 => n265_port, B2 => n11410, A => n11297, ZN 
                           => N4045);
   U17633 : OAI21_X1 port map( B1 => n264_port, B2 => n11410, A => n11301, ZN 
                           => N4046);
   U17634 : OAI21_X1 port map( B1 => n263_port, B2 => n11410, A => n11305, ZN 
                           => N4047);
   U17635 : OAI21_X1 port map( B1 => n262_port, B2 => n11410, A => n11309, ZN 
                           => N4048);
   U17636 : OAI21_X1 port map( B1 => n261_port, B2 => n11415, A => n11313, ZN 
                           => N4049);
   U17637 : OAI21_X1 port map( B1 => n260_port, B2 => n11389, A => n11317, ZN 
                           => N4050);
   U17638 : OAI21_X1 port map( B1 => n259_port, B2 => n11388, A => n11321, ZN 
                           => N4051);
   U17639 : OAI21_X1 port map( B1 => n258_port, B2 => n11388, A => n11325, ZN 
                           => N4052);
   U17640 : OAI21_X1 port map( B1 => n257_port, B2 => n11388, A => n11329, ZN 
                           => N4053);
   U17641 : OAI21_X1 port map( B1 => n256_port, B2 => n11388, A => n11077, ZN 
                           => N4055);
   U17642 : OAI21_X1 port map( B1 => n255_port, B2 => n11388, A => n11081, ZN 
                           => N4056);
   U17643 : OAI21_X1 port map( B1 => n254_port, B2 => n11388, A => n11085, ZN 
                           => N4057);
   U17644 : OAI21_X1 port map( B1 => n253_port, B2 => n11388, A => n11089, ZN 
                           => N4058);
   U17645 : OAI21_X1 port map( B1 => n252_port, B2 => n11388, A => n11093, ZN 
                           => N4059);
   U17646 : OAI21_X1 port map( B1 => n251_port, B2 => n11388, A => n11097, ZN 
                           => N4060);
   U17647 : OAI21_X1 port map( B1 => n250_port, B2 => n11388, A => n11101, ZN 
                           => N4061);
   U17648 : OAI21_X1 port map( B1 => n249_port, B2 => n11388, A => n11105, ZN 
                           => N4062);
   U17649 : OAI21_X1 port map( B1 => n248_port, B2 => n11388, A => n11109, ZN 
                           => N4063);
   U17650 : OAI21_X1 port map( B1 => n247_port, B2 => n11387, A => n11113, ZN 
                           => N4064);
   U17651 : OAI21_X1 port map( B1 => n246_port, B2 => n11387, A => n11117, ZN 
                           => N4065);
   U17652 : OAI21_X1 port map( B1 => n245_port, B2 => n11387, A => n11121, ZN 
                           => N4066);
   U17653 : OAI21_X1 port map( B1 => n244_port, B2 => n11387, A => n11125, ZN 
                           => N4067);
   U17654 : OAI21_X1 port map( B1 => n243_port, B2 => n11387, A => n11129, ZN 
                           => N4068);
   U17655 : OAI21_X1 port map( B1 => n242_port, B2 => n11387, A => n11133, ZN 
                           => N4069);
   U17656 : OAI21_X1 port map( B1 => n241_port, B2 => n11387, A => n11137, ZN 
                           => N4070);
   U17657 : OAI21_X1 port map( B1 => n240_port, B2 => n11387, A => n11141, ZN 
                           => N4071);
   U17658 : OAI21_X1 port map( B1 => n239_port, B2 => n11387, A => n11145, ZN 
                           => N4072);
   U17659 : OAI21_X1 port map( B1 => n238_port, B2 => n11387, A => n11149, ZN 
                           => N4073);
   U17660 : OAI21_X1 port map( B1 => n237_port, B2 => n11387, A => n11153, ZN 
                           => N4074);
   U17661 : OAI21_X1 port map( B1 => n236_port, B2 => n11387, A => n11157, ZN 
                           => N4075);
   U17662 : OAI21_X1 port map( B1 => n235_port, B2 => n11386, A => n11161, ZN 
                           => N4076);
   U17663 : OAI21_X1 port map( B1 => n234_port, B2 => n11386, A => n11165, ZN 
                           => N4077);
   U17664 : OAI21_X1 port map( B1 => n233_port, B2 => n11386, A => n11169, ZN 
                           => N4078);
   U17665 : OAI21_X1 port map( B1 => n232_port, B2 => n11386, A => n11173, ZN 
                           => N4079);
   U17666 : OAI21_X1 port map( B1 => n231_port, B2 => n11386, A => n11177, ZN 
                           => N4080);
   U17667 : OAI21_X1 port map( B1 => n230_port, B2 => n11386, A => n11181, ZN 
                           => N4081);
   U17668 : OAI21_X1 port map( B1 => n229_port, B2 => n11386, A => n11185, ZN 
                           => N4082);
   U17669 : OAI21_X1 port map( B1 => n228_port, B2 => n11386, A => n11189, ZN 
                           => N4083);
   U17670 : OAI21_X1 port map( B1 => n227_port, B2 => n11386, A => n11193, ZN 
                           => N4084);
   U17671 : OAI21_X1 port map( B1 => n226_port, B2 => n11386, A => n11197, ZN 
                           => N4085);
   U17672 : OAI21_X1 port map( B1 => n225_port, B2 => n11386, A => n11201, ZN 
                           => N4086);
   U17673 : OAI21_X1 port map( B1 => n224_port, B2 => n11386, A => n11205, ZN 
                           => N4087);
   U17674 : OAI21_X1 port map( B1 => n223_port, B2 => n11385, A => n11209, ZN 
                           => N4088);
   U17675 : OAI21_X1 port map( B1 => n222_port, B2 => n11385, A => n11213, ZN 
                           => N4089);
   U17676 : OAI21_X1 port map( B1 => n221_port, B2 => n11385, A => n11217, ZN 
                           => N4090);
   U17677 : OAI21_X1 port map( B1 => n220_port, B2 => n11385, A => n11221, ZN 
                           => N4091);
   U17678 : OAI21_X1 port map( B1 => n219_port, B2 => n11385, A => n11225, ZN 
                           => N4092);
   U17679 : OAI21_X1 port map( B1 => n218_port, B2 => n11385, A => n11229, ZN 
                           => N4093);
   U17680 : OAI21_X1 port map( B1 => n217_port, B2 => n11385, A => n11233, ZN 
                           => N4094);
   U17681 : OAI21_X1 port map( B1 => n216_port, B2 => n11385, A => n11237, ZN 
                           => N4095);
   U17682 : OAI21_X1 port map( B1 => n215_port, B2 => n11385, A => n11241, ZN 
                           => N4096);
   U17683 : OAI21_X1 port map( B1 => n214_port, B2 => n11385, A => n11245, ZN 
                           => N4097);
   U17684 : OAI21_X1 port map( B1 => n213_port, B2 => n11385, A => n11249, ZN 
                           => N4098);
   U17685 : OAI21_X1 port map( B1 => n212_port, B2 => n11385, A => n11253, ZN 
                           => N4099);
   U17686 : OAI21_X1 port map( B1 => n211_port, B2 => n11384, A => n11257, ZN 
                           => N4100);
   U17687 : OAI21_X1 port map( B1 => n210_port, B2 => n11384, A => n11261, ZN 
                           => N4101);
   U17688 : OAI21_X1 port map( B1 => n209_port, B2 => n11384, A => n11265, ZN 
                           => N4102);
   U17689 : OAI21_X1 port map( B1 => n208_port, B2 => n11384, A => n11269, ZN 
                           => N4103);
   U17690 : OAI21_X1 port map( B1 => n207_port, B2 => n11384, A => n11273, ZN 
                           => N4104);
   U17691 : OAI21_X1 port map( B1 => n206_port, B2 => n11384, A => n11277, ZN 
                           => N4105);
   U17692 : OAI21_X1 port map( B1 => n205_port, B2 => n11384, A => n11281, ZN 
                           => N4106);
   U17693 : OAI21_X1 port map( B1 => n204_port, B2 => n11384, A => n11285, ZN 
                           => N4107);
   U17694 : OAI21_X1 port map( B1 => n203_port, B2 => n11384, A => n11289, ZN 
                           => N4108);
   U17695 : OAI21_X1 port map( B1 => n202_port, B2 => n11384, A => n11293, ZN 
                           => N4109);
   U17696 : OAI21_X1 port map( B1 => n201_port, B2 => n11384, A => n11297, ZN 
                           => N4110);
   U17697 : OAI21_X1 port map( B1 => n200_port, B2 => n11384, A => n11301, ZN 
                           => N4111);
   U17698 : OAI21_X1 port map( B1 => n199_port, B2 => n11383, A => n11305, ZN 
                           => N4112);
   U17699 : OAI21_X1 port map( B1 => n198_port, B2 => n11383, A => n11309, ZN 
                           => N4113);
   U17700 : OAI21_X1 port map( B1 => n197_port, B2 => n11383, A => n11313, ZN 
                           => N4114);
   U17701 : OAI21_X1 port map( B1 => n196_port, B2 => n11383, A => n11317, ZN 
                           => N4115);
   U17702 : OAI21_X1 port map( B1 => n195_port, B2 => n11383, A => n11321, ZN 
                           => N4116);
   U17703 : OAI21_X1 port map( B1 => n194_port, B2 => n11383, A => n11325, ZN 
                           => N4117);
   U17704 : OAI21_X1 port map( B1 => n193_port, B2 => n11383, A => n11329, ZN 
                           => N4118);
   U17705 : OAI21_X1 port map( B1 => n192_port, B2 => n11383, A => n11077, ZN 
                           => N4120);
   U17706 : OAI21_X1 port map( B1 => n191_port, B2 => n11383, A => n11081, ZN 
                           => N4121);
   U17707 : OAI21_X1 port map( B1 => n190_port, B2 => n11383, A => n11085, ZN 
                           => N4122);
   U17708 : OAI21_X1 port map( B1 => n189_port, B2 => n11383, A => n11089, ZN 
                           => N4123);
   U17709 : OAI21_X1 port map( B1 => n188_port, B2 => n11382, A => n11093, ZN 
                           => N4124);
   U17710 : OAI21_X1 port map( B1 => n187_port, B2 => n11382, A => n11097, ZN 
                           => N4125);
   U17711 : OAI21_X1 port map( B1 => n186_port, B2 => n11382, A => n11101, ZN 
                           => N4126);
   U17712 : OAI21_X1 port map( B1 => n185_port, B2 => n11382, A => n11105, ZN 
                           => N4127);
   U17713 : OAI21_X1 port map( B1 => n184_port, B2 => n11382, A => n11109, ZN 
                           => N4128);
   U17714 : OAI21_X1 port map( B1 => n183_port, B2 => n11382, A => n11113, ZN 
                           => N4129);
   U17715 : OAI21_X1 port map( B1 => n182_port, B2 => n11382, A => n11117, ZN 
                           => N4130);
   U17716 : OAI21_X1 port map( B1 => n181_port, B2 => n11382, A => n11121, ZN 
                           => N4131);
   U17717 : OAI21_X1 port map( B1 => n180_port, B2 => n11382, A => n11125, ZN 
                           => N4132);
   U17718 : OAI21_X1 port map( B1 => n179_port, B2 => n11382, A => n11129, ZN 
                           => N4133);
   U17719 : OAI21_X1 port map( B1 => n178_port, B2 => n11382, A => n11133, ZN 
                           => N4134);
   U17720 : OAI21_X1 port map( B1 => n177_port, B2 => n11382, A => n11137, ZN 
                           => N4135);
   U17721 : OAI21_X1 port map( B1 => n176_port, B2 => n11381, A => n11141, ZN 
                           => N4136);
   U17722 : OAI21_X1 port map( B1 => n175_port, B2 => n11381, A => n11145, ZN 
                           => N4137);
   U17723 : OAI21_X1 port map( B1 => n174_port, B2 => n11381, A => n11149, ZN 
                           => N4138);
   U17724 : OAI21_X1 port map( B1 => n173_port, B2 => n11381, A => n11153, ZN 
                           => N4139);
   U17725 : OAI21_X1 port map( B1 => n172_port, B2 => n11381, A => n11157, ZN 
                           => N4140);
   U17726 : OAI21_X1 port map( B1 => n171_port, B2 => n11381, A => n11161, ZN 
                           => N4141);
   U17727 : OAI21_X1 port map( B1 => n170_port, B2 => n11381, A => n11165, ZN 
                           => N4142);
   U17728 : OAI21_X1 port map( B1 => n169_port, B2 => n11381, A => n11169, ZN 
                           => N4143);
   U17729 : OAI21_X1 port map( B1 => n168_port, B2 => n11381, A => n11173, ZN 
                           => N4144);
   U17730 : OAI21_X1 port map( B1 => n167_port, B2 => n11381, A => n11177, ZN 
                           => N4145);
   U17731 : OAI21_X1 port map( B1 => n166_port, B2 => n11381, A => n11181, ZN 
                           => N4146);
   U17732 : OAI21_X1 port map( B1 => n165_port, B2 => n11381, A => n11185, ZN 
                           => N4147);
   U17733 : OAI21_X1 port map( B1 => n164_port, B2 => n11380, A => n11189, ZN 
                           => N4148);
   U17734 : OAI21_X1 port map( B1 => n163_port, B2 => n11380, A => n11193, ZN 
                           => N4149);
   U17735 : OAI21_X1 port map( B1 => n162_port, B2 => n11380, A => n11197, ZN 
                           => N4150);
   U17736 : OAI21_X1 port map( B1 => n161_port, B2 => n11380, A => n11201, ZN 
                           => N4151);
   U17737 : OAI21_X1 port map( B1 => n160_port, B2 => n11380, A => n11205, ZN 
                           => N4152);
   U17738 : OAI21_X1 port map( B1 => n159_port, B2 => n11380, A => n11209, ZN 
                           => N4153);
   U17739 : OAI21_X1 port map( B1 => n158_port, B2 => n11380, A => n11213, ZN 
                           => N4154);
   U17740 : OAI21_X1 port map( B1 => n157_port, B2 => n11380, A => n11217, ZN 
                           => N4155);
   U17741 : OAI21_X1 port map( B1 => n156_port, B2 => n11380, A => n11221, ZN 
                           => N4156);
   U17742 : OAI21_X1 port map( B1 => n155_port, B2 => n11380, A => n11225, ZN 
                           => N4157);
   U17743 : OAI21_X1 port map( B1 => n154_port, B2 => n11380, A => n11229, ZN 
                           => N4158);
   U17744 : OAI21_X1 port map( B1 => n153_port, B2 => n11380, A => n11233, ZN 
                           => N4159);
   U17745 : OAI21_X1 port map( B1 => n152_port, B2 => n11379, A => n11237, ZN 
                           => N4160);
   U17746 : OAI21_X1 port map( B1 => n151_port, B2 => n11379, A => n11241, ZN 
                           => N4161);
   U17747 : OAI21_X1 port map( B1 => n150_port, B2 => n11379, A => n11245, ZN 
                           => N4162);
   U17748 : OAI21_X1 port map( B1 => n149_port, B2 => n11379, A => n11249, ZN 
                           => N4163);
   U17749 : OAI21_X1 port map( B1 => n148_port, B2 => n11379, A => n11253, ZN 
                           => N4164);
   U17750 : OAI21_X1 port map( B1 => n147_port, B2 => n11379, A => n11257, ZN 
                           => N4165);
   U17751 : OAI21_X1 port map( B1 => n146_port, B2 => n11379, A => n11261, ZN 
                           => N4166);
   U17752 : OAI21_X1 port map( B1 => n145_port, B2 => n11379, A => n11265, ZN 
                           => N4167);
   U17753 : OAI21_X1 port map( B1 => n144_port, B2 => n11379, A => n11269, ZN 
                           => N4168);
   U17754 : OAI21_X1 port map( B1 => n143_port, B2 => n11379, A => n11273, ZN 
                           => N4169);
   U17755 : OAI21_X1 port map( B1 => n142_port, B2 => n11379, A => n11277, ZN 
                           => N4170);
   U17756 : OAI21_X1 port map( B1 => n141_port, B2 => n11379, A => n11281, ZN 
                           => N4171);
   U17757 : OAI21_X1 port map( B1 => n140_port, B2 => n11378, A => n11285, ZN 
                           => N4172);
   U17758 : OAI21_X1 port map( B1 => n139_port, B2 => n11378, A => n11289, ZN 
                           => N4173);
   U17759 : OAI21_X1 port map( B1 => n138_port, B2 => n11378, A => n11293, ZN 
                           => N4174);
   U17760 : OAI21_X1 port map( B1 => n137_port, B2 => n11378, A => n11297, ZN 
                           => N4175);
   U17761 : OAI21_X1 port map( B1 => n136_port, B2 => n11378, A => n11301, ZN 
                           => N4176);
   U17762 : OAI21_X1 port map( B1 => n135_port, B2 => n11378, A => n11305, ZN 
                           => N4177);
   U17763 : OAI21_X1 port map( B1 => n134_port, B2 => n11378, A => n11309, ZN 
                           => N4178);
   U17764 : OAI21_X1 port map( B1 => n133_port, B2 => n11378, A => n11313, ZN 
                           => N4179);
   U17765 : OAI21_X1 port map( B1 => n132_port, B2 => n11383, A => n11317, ZN 
                           => N4180);
   U17766 : OAI21_X1 port map( B1 => n131_port, B2 => n11399, A => n11321, ZN 
                           => N4181);
   U17767 : OAI21_X1 port map( B1 => n130_port, B2 => n11399, A => n11325, ZN 
                           => N4182);
   U17768 : OAI21_X1 port map( B1 => n129_port, B2 => n11399, A => n11329, ZN 
                           => N4183);
   U17769 : OAI21_X1 port map( B1 => n128_port, B2 => n11399, A => n11077, ZN 
                           => N4185);
   U17770 : OAI21_X1 port map( B1 => n127_port, B2 => n11399, A => n11081, ZN 
                           => N4186);
   U17771 : OAI21_X1 port map( B1 => n126_port, B2 => n11399, A => n11085, ZN 
                           => N4187);
   U17772 : OAI21_X1 port map( B1 => n125_port, B2 => n11399, A => n11089, ZN 
                           => N4188);
   U17773 : OAI21_X1 port map( B1 => n124_port, B2 => n11399, A => n11093, ZN 
                           => N4189);
   U17774 : OAI21_X1 port map( B1 => n123_port, B2 => n11399, A => n11097, ZN 
                           => N4190);
   U17775 : OAI21_X1 port map( B1 => n122_port, B2 => n11398, A => n11101, ZN 
                           => N4191);
   U17776 : OAI21_X1 port map( B1 => n121_port, B2 => n11398, A => n11105, ZN 
                           => N4192);
   U17777 : OAI21_X1 port map( B1 => n120_port, B2 => n11398, A => n11109, ZN 
                           => N4193);
   U17778 : OAI21_X1 port map( B1 => n119_port, B2 => n11398, A => n11113, ZN 
                           => N4194);
   U17779 : OAI21_X1 port map( B1 => n118_port, B2 => n11398, A => n11117, ZN 
                           => N4195);
   U17780 : OAI21_X1 port map( B1 => n117_port, B2 => n11398, A => n11121, ZN 
                           => N4196);
   U17781 : OAI21_X1 port map( B1 => n116_port, B2 => n11398, A => n11125, ZN 
                           => N4197);
   U17782 : OAI21_X1 port map( B1 => n115_port, B2 => n11398, A => n11129, ZN 
                           => N4198);
   U17783 : OAI21_X1 port map( B1 => n114_port, B2 => n11398, A => n11133, ZN 
                           => N4199);
   U17784 : OAI21_X1 port map( B1 => n113_port, B2 => n11398, A => n11137, ZN 
                           => N4200);
   U17785 : OAI21_X1 port map( B1 => n112_port, B2 => n11398, A => n11141, ZN 
                           => N4201);
   U17786 : OAI21_X1 port map( B1 => n111_port, B2 => n11398, A => n11145, ZN 
                           => N4202);
   U17787 : OAI21_X1 port map( B1 => n110_port, B2 => n11397, A => n11149, ZN 
                           => N4203);
   U17788 : OAI21_X1 port map( B1 => n109_port, B2 => n11397, A => n11153, ZN 
                           => N4204);
   U17789 : OAI21_X1 port map( B1 => n108_port, B2 => n11397, A => n11157, ZN 
                           => N4205);
   U17790 : OAI21_X1 port map( B1 => n107_port, B2 => n11397, A => n11161, ZN 
                           => N4206);
   U17791 : OAI21_X1 port map( B1 => n106_port, B2 => n11397, A => n11165, ZN 
                           => N4207);
   U17792 : OAI21_X1 port map( B1 => n105_port, B2 => n11397, A => n11169, ZN 
                           => N4208);
   U17793 : OAI21_X1 port map( B1 => n104_port, B2 => n11397, A => n11173, ZN 
                           => N4209);
   U17794 : OAI21_X1 port map( B1 => n103_port, B2 => n11397, A => n11177, ZN 
                           => N4210);
   U17795 : OAI21_X1 port map( B1 => n102_port, B2 => n11397, A => n11181, ZN 
                           => N4211);
   U17796 : OAI21_X1 port map( B1 => n101_port, B2 => n11397, A => n11185, ZN 
                           => N4212);
   U17797 : OAI21_X1 port map( B1 => n100_port, B2 => n11397, A => n11189, ZN 
                           => N4213);
   U17798 : OAI21_X1 port map( B1 => n99_port, B2 => n11397, A => n11193, ZN =>
                           N4214);
   U17799 : OAI21_X1 port map( B1 => n98_port, B2 => n11396, A => n11197, ZN =>
                           N4215);
   U17800 : OAI21_X1 port map( B1 => n97_port, B2 => n11396, A => n11201, ZN =>
                           N4216);
   U17801 : OAI21_X1 port map( B1 => n96_port, B2 => n11396, A => n11205, ZN =>
                           N4217);
   U17802 : OAI21_X1 port map( B1 => n95_port, B2 => n11396, A => n11209, ZN =>
                           N4218);
   U17803 : OAI21_X1 port map( B1 => n94_port, B2 => n11396, A => n11213, ZN =>
                           N4219);
   U17804 : OAI21_X1 port map( B1 => n93_port, B2 => n11396, A => n11217, ZN =>
                           N4220);
   U17805 : OAI21_X1 port map( B1 => n92_port, B2 => n11396, A => n11221, ZN =>
                           N4221);
   U17806 : OAI21_X1 port map( B1 => n91_port, B2 => n11396, A => n11225, ZN =>
                           N4222);
   U17807 : OAI21_X1 port map( B1 => n90_port, B2 => n11396, A => n11229, ZN =>
                           N4223);
   U17808 : OAI21_X1 port map( B1 => n89_port, B2 => n11396, A => n11233, ZN =>
                           N4224);
   U17809 : OAI21_X1 port map( B1 => n88_port, B2 => n11396, A => n11237, ZN =>
                           N4225);
   U17810 : OAI21_X1 port map( B1 => n87_port, B2 => n11396, A => n11241, ZN =>
                           N4226);
   U17811 : OAI21_X1 port map( B1 => n86_port, B2 => n11395, A => n11245, ZN =>
                           N4227);
   U17812 : OAI21_X1 port map( B1 => n85_port, B2 => n11395, A => n11249, ZN =>
                           N4228);
   U17813 : OAI21_X1 port map( B1 => n84_port, B2 => n11395, A => n11253, ZN =>
                           N4229);
   U17814 : OAI21_X1 port map( B1 => n83_port, B2 => n11395, A => n11257, ZN =>
                           N4230);
   U17815 : OAI21_X1 port map( B1 => n82_port, B2 => n11395, A => n11261, ZN =>
                           N4231);
   U17816 : OAI21_X1 port map( B1 => n81_port, B2 => n11395, A => n11265, ZN =>
                           N4232);
   U17817 : OAI21_X1 port map( B1 => n80_port, B2 => n11395, A => n11269, ZN =>
                           N4233);
   U17818 : OAI21_X1 port map( B1 => n79_port, B2 => n11395, A => n11273, ZN =>
                           N4234);
   U17819 : OAI21_X1 port map( B1 => n78_port, B2 => n11395, A => n11277, ZN =>
                           N4235);
   U17820 : OAI21_X1 port map( B1 => n77_port, B2 => n11395, A => n11281, ZN =>
                           N4236);
   U17821 : OAI21_X1 port map( B1 => n76_port, B2 => n11395, A => n11285, ZN =>
                           N4237);
   U17822 : OAI21_X1 port map( B1 => n75_port, B2 => n11395, A => n11289, ZN =>
                           N4238);
   U17823 : OAI21_X1 port map( B1 => n74_port, B2 => n11394, A => n11293, ZN =>
                           N4239);
   U17824 : OAI21_X1 port map( B1 => n73_port, B2 => n11394, A => n11297, ZN =>
                           N4240);
   U17825 : OAI21_X1 port map( B1 => n72_port, B2 => n11394, A => n11301, ZN =>
                           N4241);
   U17826 : OAI21_X1 port map( B1 => n71_port, B2 => n11394, A => n11305, ZN =>
                           N4242);
   U17827 : OAI21_X1 port map( B1 => n70_port, B2 => n11394, A => n11309, ZN =>
                           N4243);
   U17828 : OAI21_X1 port map( B1 => n69_port, B2 => n11394, A => n11313, ZN =>
                           N4244);
   U17829 : OAI21_X1 port map( B1 => n68_port, B2 => n11394, A => n11317, ZN =>
                           N4245);
   U17830 : OAI21_X1 port map( B1 => n67_port, B2 => n11394, A => n11321, ZN =>
                           N4246);
   U17831 : OAI21_X1 port map( B1 => n66_port, B2 => n11394, A => n11325, ZN =>
                           N4247);
   U17832 : OAI21_X1 port map( B1 => n65_port, B2 => n11394, A => n11329, ZN =>
                           N4248);
   U17833 : OAI21_X1 port map( B1 => n64_port, B2 => n11394, A => n11077, ZN =>
                           N4250);
   U17834 : OAI21_X1 port map( B1 => n63_port, B2 => n11393, A => n11081, ZN =>
                           N4251);
   U17835 : OAI21_X1 port map( B1 => n62_port, B2 => n11393, A => n11085, ZN =>
                           N4252);
   U17836 : OAI21_X1 port map( B1 => n61_port, B2 => n11393, A => n11089, ZN =>
                           N4253);
   U17837 : OAI21_X1 port map( B1 => n60_port, B2 => n11393, A => n11093, ZN =>
                           N4254);
   U17838 : OAI21_X1 port map( B1 => n59_port, B2 => n11393, A => n11097, ZN =>
                           N4255);
   U17839 : OAI21_X1 port map( B1 => n58_port, B2 => n11393, A => n11101, ZN =>
                           N4256);
   U17840 : OAI21_X1 port map( B1 => n57_port, B2 => n11393, A => n11105, ZN =>
                           N4257);
   U17841 : OAI21_X1 port map( B1 => n56_port, B2 => n11393, A => n11109, ZN =>
                           N4258);
   U17842 : OAI21_X1 port map( B1 => n55_port, B2 => n11393, A => n11113, ZN =>
                           N4259);
   U17843 : OAI21_X1 port map( B1 => n54_port, B2 => n11393, A => n11117, ZN =>
                           N4260);
   U17844 : OAI21_X1 port map( B1 => n53_port, B2 => n11393, A => n11121, ZN =>
                           N4261);
   U17845 : OAI21_X1 port map( B1 => n52_port, B2 => n11393, A => n11125, ZN =>
                           N4262);
   U17846 : OAI21_X1 port map( B1 => n51_port, B2 => n11392, A => n11129, ZN =>
                           N4263);
   U17847 : OAI21_X1 port map( B1 => n50_port, B2 => n11392, A => n11133, ZN =>
                           N4264);
   U17848 : OAI21_X1 port map( B1 => n49_port, B2 => n11392, A => n11137, ZN =>
                           N4265);
   U17849 : OAI21_X1 port map( B1 => n48_port, B2 => n11392, A => n11141, ZN =>
                           N4266);
   U17850 : OAI21_X1 port map( B1 => n47_port, B2 => n11392, A => n11145, ZN =>
                           N4267);
   U17851 : OAI21_X1 port map( B1 => n46_port, B2 => n11392, A => n11149, ZN =>
                           N4268);
   U17852 : OAI21_X1 port map( B1 => n45_port, B2 => n11392, A => n11153, ZN =>
                           N4269);
   U17853 : OAI21_X1 port map( B1 => n44_port, B2 => n11392, A => n11157, ZN =>
                           N4270);
   U17854 : OAI21_X1 port map( B1 => n43_port, B2 => n11392, A => n11161, ZN =>
                           N4271);
   U17855 : OAI21_X1 port map( B1 => n42_port, B2 => n11392, A => n11165, ZN =>
                           N4272);
   U17856 : OAI21_X1 port map( B1 => n41_port, B2 => n11392, A => n11169, ZN =>
                           N4273);
   U17857 : OAI21_X1 port map( B1 => n40_port, B2 => n11392, A => n11173, ZN =>
                           N4274);
   U17858 : OAI21_X1 port map( B1 => n39_port, B2 => n11391, A => n11177, ZN =>
                           N4275);
   U17859 : OAI21_X1 port map( B1 => n38_port, B2 => n11391, A => n11181, ZN =>
                           N4276);
   U17860 : OAI21_X1 port map( B1 => n37_port, B2 => n11391, A => n11185, ZN =>
                           N4277);
   U17861 : OAI21_X1 port map( B1 => n36_port, B2 => n11391, A => n11189, ZN =>
                           N4278);
   U17862 : OAI21_X1 port map( B1 => n35_port, B2 => n11391, A => n11193, ZN =>
                           N4279);
   U17863 : OAI21_X1 port map( B1 => n34_port, B2 => n11391, A => n11197, ZN =>
                           N4280);
   U17864 : OAI21_X1 port map( B1 => n33_port, B2 => n11391, A => n11201, ZN =>
                           N4281);
   U17865 : OAI21_X1 port map( B1 => n32_port, B2 => n11391, A => n11205, ZN =>
                           N4282);
   U17866 : OAI21_X1 port map( B1 => n31_port, B2 => n11391, A => n11209, ZN =>
                           N4283);
   U17867 : OAI21_X1 port map( B1 => n30_port, B2 => n11391, A => n11213, ZN =>
                           N4284);
   U17868 : OAI21_X1 port map( B1 => n29_port, B2 => n11391, A => n11217, ZN =>
                           N4285);
   U17869 : OAI21_X1 port map( B1 => n28_port, B2 => n11391, A => n11221, ZN =>
                           N4286);
   U17870 : OAI21_X1 port map( B1 => n27_port, B2 => n11390, A => n11225, ZN =>
                           N4287);
   U17871 : OAI21_X1 port map( B1 => n26_port, B2 => n11390, A => n11229, ZN =>
                           N4288);
   U17872 : OAI21_X1 port map( B1 => n25_port, B2 => n11390, A => n11233, ZN =>
                           N4289);
   U17873 : OAI21_X1 port map( B1 => n24_port, B2 => n11390, A => n11237, ZN =>
                           N4290);
   U17874 : OAI21_X1 port map( B1 => n23_port, B2 => n11390, A => n11241, ZN =>
                           N4291);
   U17875 : OAI21_X1 port map( B1 => n22_port, B2 => n11390, A => n11245, ZN =>
                           N4292);
   U17876 : OAI21_X1 port map( B1 => n21, B2 => n11390, A => n11249, ZN => 
                           N4293);
   U17877 : OAI21_X1 port map( B1 => n20, B2 => n11390, A => n11253, ZN => 
                           N4294);
   U17878 : OAI21_X1 port map( B1 => n19, B2 => n11390, A => n11257, ZN => 
                           N4295);
   U17879 : OAI21_X1 port map( B1 => n18, B2 => n11390, A => n11261, ZN => 
                           N4296);
   U17880 : OAI21_X1 port map( B1 => n17, B2 => n11390, A => n11265, ZN => 
                           N4297);
   U17881 : OAI21_X1 port map( B1 => n16, B2 => n11390, A => n11269, ZN => 
                           N4298);
   U17882 : OAI21_X1 port map( B1 => n15, B2 => n11389, A => n11273, ZN => 
                           N4299);
   U17883 : OAI21_X1 port map( B1 => n14, B2 => n11389, A => n11277, ZN => 
                           N4300);
   U17884 : OAI21_X1 port map( B1 => n13, B2 => n11389, A => n11281, ZN => 
                           N4301);
   U17885 : OAI21_X1 port map( B1 => n12, B2 => n11389, A => n11285, ZN => 
                           N4302);
   U17886 : OAI21_X1 port map( B1 => n11, B2 => n11389, A => n11289, ZN => 
                           N4303);
   U17887 : OAI21_X1 port map( B1 => n10, B2 => n11389, A => n11293, ZN => 
                           N4304);
   U17888 : OAI21_X1 port map( B1 => n9, B2 => n11389, A => n11297, ZN => N4305
                           );
   U17889 : OAI21_X1 port map( B1 => n8, B2 => n11389, A => n11301, ZN => N4306
                           );
   U17890 : OAI21_X1 port map( B1 => n7, B2 => n11389, A => n11305, ZN => N4307
                           );
   U17891 : OAI21_X1 port map( B1 => n6, B2 => n11389, A => n11309, ZN => N4308
                           );
   U17892 : OAI21_X1 port map( B1 => n5, B2 => n11389, A => n11313, ZN => N4309
                           );
   U17893 : OAI21_X1 port map( B1 => n4, B2 => n11394, A => n11317, ZN => N4310
                           );
   U17894 : OAI21_X1 port map( B1 => n3, B2 => n11399, A => n11321, ZN => N4311
                           );
   U17895 : OAI21_X1 port map( B1 => n2, B2 => n11340, A => n11325, ZN => N4312
                           );
   U17896 : OAI21_X1 port map( B1 => n1, B2 => n11421, A => n11329, ZN => N4313
                           );
   U17897 : OAI21_X1 port map( B1 => n678_port, B2 => n11335, A => n11180, ZN 
                           => N3626);
   U17898 : OAI21_X1 port map( B1 => n677_port, B2 => n11335, A => n11184, ZN 
                           => N3627);
   U17899 : OAI21_X1 port map( B1 => n675_port, B2 => n11335, A => n11192, ZN 
                           => N3629);
   U17900 : OAI21_X1 port map( B1 => n674_port, B2 => n11335, A => n11196, ZN 
                           => N3630);
   U17901 : OAI21_X1 port map( B1 => n671_port, B2 => n11335, A => n11208, ZN 
                           => N3633);
   U17902 : OAI21_X1 port map( B1 => n669_port, B2 => n11335, A => n11216, ZN 
                           => N3635);
   U17903 : OAI21_X1 port map( B1 => n667_port, B2 => n11335, A => n11224, ZN 
                           => N3637);
   U17904 : OAI21_X1 port map( B1 => n663_port, B2 => n11335, A => n11240, ZN 
                           => N3641);
   U17905 : INV_X1 port map( A => ADD_WR(2), ZN => n6229);
   U17906 : INV_X1 port map( A => ADD_WR(0), ZN => n6231);
   U17907 : INV_X1 port map( A => ADD_WR(1), ZN => n6230);
   U17908 : INV_X1 port map( A => ADD_WR(3), ZN => n6228);
   U17909 : INV_X1 port map( A => ADD_RD2(3), ZN => n6242);
   U17910 : INV_X1 port map( A => ADD_RD1(3), ZN => n6233);
   U17911 : BUF_X1 port map( A => n7301, Z => n11011);
   U17912 : NOR3_X1 port map( A1 => n6249, A2 => ADD_RD2(1), A3 => n6247, ZN =>
                           n7301);
   U17913 : BUF_X1 port map( A => n7298, Z => n11046);
   U17914 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n7298);
   U17915 : BUF_X1 port map( A => n8481, Z => n10786);
   U17916 : NOR3_X1 port map( A1 => n6240, A2 => ADD_RD1(1), A3 => n6238, ZN =>
                           n8481);
   U17917 : BUF_X1 port map( A => n8478, Z => n10821);
   U17918 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n8478);
   U17919 : BUF_X1 port map( A => n7297, Z => n11064);
   U17920 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n6248, 
                           ZN => n7297);
   U17921 : BUF_X1 port map( A => n8477, Z => n10839);
   U17922 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n6239, 
                           ZN => n8477);
   U17923 : INV_X1 port map( A => ADD_WR(4), ZN => n6227);
   U17924 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n11335, ZN => n7274);
   U17925 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n11334, ZN => n7273);
   U17926 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n11335, ZN => n7272);
   U17927 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n11334, ZN => n7271);
   U17928 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n11334, ZN => n7270);
   U17929 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n11335, ZN => n7269);
   U17930 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n11335, ZN => n7268);
   U17931 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n11334, ZN => n7267);
   U17932 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n11334, ZN => n7266);
   U17933 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n11334, ZN => n7265);
   U17934 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n11333, ZN => n7264);
   U17935 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n11334, ZN => n7263);
   U17936 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n11334, ZN => n7262);
   U17937 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n11334, ZN => n7261);
   U17938 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n11334, ZN => n7260);
   U17939 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n11334, ZN => n7259);
   U17940 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n11333, ZN => n7258);
   U17941 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n11333, ZN => n7257);
   U17942 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n11334, ZN => n7256);
   U17943 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n11333, ZN => n7255);
   U17944 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n11333, ZN => n7254);
   U17945 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n11333, ZN => n7253);
   U17946 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n11333, ZN => n7252);
   U17947 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n11333, ZN => n7251);
   U17948 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n11333, ZN => n7250);
   U17949 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n11333, ZN => n7249);
   U17950 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n11333, ZN => n7248);
   U17951 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n11332, ZN => n7247);
   U17952 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n11332, ZN => n7246);
   U17953 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n11332, ZN => n7245);
   U17954 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n11332, ZN => n7244);
   U17955 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n11333, ZN => n7243);
   U17956 : NAND2_X1 port map( A1 => DATAIN(32), A2 => n11332, ZN => n7242);
   U17957 : NAND2_X1 port map( A1 => DATAIN(33), A2 => n11332, ZN => n7241);
   U17958 : NAND2_X1 port map( A1 => DATAIN(34), A2 => n11332, ZN => n7240);
   U17959 : NAND2_X1 port map( A1 => DATAIN(35), A2 => n11332, ZN => n7239);
   U17960 : NAND2_X1 port map( A1 => DATAIN(36), A2 => n11332, ZN => n7238);
   U17961 : NAND2_X1 port map( A1 => DATAIN(37), A2 => n11332, ZN => n7237);
   U17962 : NAND2_X1 port map( A1 => DATAIN(38), A2 => n11332, ZN => n7236);
   U17963 : NAND2_X1 port map( A1 => DATAIN(39), A2 => n11331, ZN => n7235);
   U17964 : NAND2_X1 port map( A1 => DATAIN(40), A2 => n11331, ZN => n7234);
   U17965 : NAND2_X1 port map( A1 => DATAIN(41), A2 => n11331, ZN => n7233);
   U17966 : NAND2_X1 port map( A1 => DATAIN(42), A2 => n11331, ZN => n7232);
   U17967 : NAND2_X1 port map( A1 => DATAIN(43), A2 => n11331, ZN => n7231);
   U17968 : NAND2_X1 port map( A1 => DATAIN(44), A2 => n11331, ZN => n7230);
   U17969 : NAND2_X1 port map( A1 => DATAIN(45), A2 => n11331, ZN => n7229);
   U17970 : NAND2_X1 port map( A1 => DATAIN(46), A2 => n11331, ZN => n7228);
   U17971 : NAND2_X1 port map( A1 => DATAIN(47), A2 => n11331, ZN => n7227);
   U17972 : NAND2_X1 port map( A1 => DATAIN(48), A2 => n11331, ZN => n7226);
   U17973 : NAND2_X1 port map( A1 => DATAIN(49), A2 => n11331, ZN => n7225);
   U17974 : NAND2_X1 port map( A1 => DATAIN(50), A2 => n11331, ZN => n7224);
   U17975 : NAND2_X1 port map( A1 => DATAIN(51), A2 => n11330, ZN => n7223);
   U17976 : NAND2_X1 port map( A1 => DATAIN(52), A2 => n11330, ZN => n7222);
   U17977 : NAND2_X1 port map( A1 => DATAIN(53), A2 => n11330, ZN => n7221);
   U17978 : NAND2_X1 port map( A1 => DATAIN(54), A2 => n11330, ZN => n7220);
   U17979 : NAND2_X1 port map( A1 => DATAIN(55), A2 => n11330, ZN => n7219);
   U17980 : NAND2_X1 port map( A1 => DATAIN(56), A2 => n11330, ZN => n7218);
   U17981 : NAND2_X1 port map( A1 => DATAIN(57), A2 => n11330, ZN => n7217);
   U17982 : NAND2_X1 port map( A1 => DATAIN(58), A2 => n11330, ZN => n7216);
   U17983 : NAND2_X1 port map( A1 => DATAIN(59), A2 => n11330, ZN => n7215);
   U17984 : NAND2_X1 port map( A1 => DATAIN(60), A2 => n11330, ZN => n7214);
   U17985 : NAND2_X1 port map( A1 => DATAIN(61), A2 => n11330, ZN => n7213);
   U17986 : NAND2_X1 port map( A1 => DATAIN(62), A2 => n11330, ZN => n7212);
   U17987 : NAND2_X1 port map( A1 => DATAIN(63), A2 => n11332, ZN => n7211);
   U17988 : INV_X1 port map( A => RESET, ZN => n6226);
   U17989 : BUF_X1 port map( A => n7305, Z => n10986);
   U17990 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => n6241, ZN => n7305);
   U17991 : BUF_X1 port map( A => n8485, Z => n10761);
   U17992 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => n6232, ZN => n8485);
   U17993 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_0_port, A2 => n11766, ZN 
                           => N22);
   U17994 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_1_port, A2 => n11767, ZN 
                           => N23);
   U17995 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_2_port, A2 => n11768, ZN 
                           => N24);
   U17996 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_3_port, A2 => n11768, ZN 
                           => N25);
   U17997 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_4_port, A2 => n11769, ZN 
                           => N26);
   U17998 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_5_port, A2 => n11770, ZN 
                           => N27);
   U17999 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_6_port, A2 => n11771, ZN 
                           => N28);
   U18000 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_7_port, A2 => n11772, ZN 
                           => N29);
   U18001 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_8_port, A2 => n11773, ZN 
                           => N30);
   U18002 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_9_port, A2 => n11774, ZN 
                           => N31);
   U18003 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_10_port, A2 => n11775, ZN
                           => N32);
   U18004 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_11_port, A2 => n11776, ZN
                           => N33);
   U18005 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_12_port, A2 => n11777, ZN
                           => N34);
   U18006 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_13_port, A2 => n11778, ZN
                           => N35);
   U18007 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_14_port, A2 => n11779, ZN
                           => N36);
   U18008 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_15_port, A2 => n11779, ZN
                           => N37);
   U18009 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_16_port, A2 => n11780, ZN
                           => N38);
   U18010 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_17_port, A2 => n11781, ZN
                           => N39);
   U18011 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_18_port, A2 => n11782, ZN
                           => N40);
   U18012 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_19_port, A2 => n11783, ZN
                           => N41);
   U18013 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_20_port, A2 => n11784, ZN
                           => N42);
   U18014 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_21_port, A2 => n11785, ZN
                           => N43);
   U18015 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_22_port, A2 => n11786, ZN
                           => N44);
   U18016 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_23_port, A2 => n11787, ZN
                           => N45);
   U18017 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_24_port, A2 => n11788, ZN
                           => N46);
   U18018 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_25_port, A2 => n11789, ZN
                           => N47);
   U18019 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_26_port, A2 => n11790, ZN
                           => N48);
   U18020 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_27_port, A2 => n11790, ZN
                           => N49);
   U18021 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_28_port, A2 => n11791, ZN
                           => N50);
   U18022 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_29_port, A2 => n11792, ZN
                           => N51);
   U18023 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_30_port, A2 => n11793, ZN
                           => N52);
   U18024 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_31_port, A2 => n11794, ZN
                           => N53);
   U18025 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_32_port, A2 => n11795, ZN
                           => N54);
   U18026 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_33_port, A2 => n11796, ZN
                           => N55);
   U18027 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_34_port, A2 => n11797, ZN
                           => N56);
   U18028 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_35_port, A2 => n11798, ZN
                           => N57);
   U18029 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_36_port, A2 => n11799, ZN
                           => N58);
   U18030 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_37_port, A2 => n11800, ZN
                           => N59);
   U18031 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_38_port, A2 => n11801, ZN
                           => N60);
   U18032 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_39_port, A2 => n11801, ZN
                           => N61);
   U18033 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_40_port, A2 => n11802, ZN
                           => N62);
   U18034 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_41_port, A2 => n11803, ZN
                           => N63);
   U18035 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_42_port, A2 => n11804, ZN
                           => N64);
   U18036 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_43_port, A2 => n11805, ZN
                           => N65);
   U18037 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_44_port, A2 => n11806, ZN
                           => N66);
   U18038 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_45_port, A2 => n11807, ZN
                           => N67);
   U18039 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_46_port, A2 => n11808, ZN
                           => N68);
   U18040 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_47_port, A2 => n11809, ZN
                           => N69);
   U18041 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_48_port, A2 => n11810, ZN
                           => N70);
   U18042 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_49_port, A2 => n11811, ZN
                           => N71);
   U18043 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_50_port, A2 => n11812, ZN
                           => N72);
   U18044 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_51_port, A2 => n11812, ZN
                           => N73);
   U18045 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_52_port, A2 => n11813, ZN
                           => N74);
   U18046 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_53_port, A2 => n11814, ZN
                           => N75);
   U18047 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_54_port, A2 => n11815, ZN
                           => N76);
   U18048 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_55_port, A2 => n11816, ZN
                           => N77);
   U18049 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_56_port, A2 => n11817, ZN
                           => N78);
   U18050 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_57_port, A2 => n11818, ZN
                           => N79);
   U18051 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_58_port, A2 => n11819, ZN
                           => N80);
   U18052 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_59_port, A2 => n11820, ZN
                           => N81);
   U18053 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_60_port, A2 => n11821, ZN
                           => N82);
   U18054 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_61_port, A2 => n11822, ZN
                           => N83);
   U18055 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_62_port, A2 => n11823, ZN
                           => N84);
   U18056 : AND2_X1 port map( A1 => NEXT_REGISTERS_31_63_port, A2 => n11823, ZN
                           => N85);
   U18057 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_0_port, A2 => n11824, ZN 
                           => N86);
   U18058 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_1_port, A2 => n11825, ZN 
                           => N87);
   U18059 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_2_port, A2 => n11826, ZN 
                           => N88);
   U18060 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_3_port, A2 => n11827, ZN 
                           => N89);
   U18061 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_4_port, A2 => n11828, ZN 
                           => N90);
   U18062 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_5_port, A2 => n11829, ZN 
                           => N91);
   U18063 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_6_port, A2 => n11830, ZN 
                           => N92);
   U18064 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_7_port, A2 => n11831, ZN 
                           => N93);
   U18065 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_8_port, A2 => n11832, ZN 
                           => N94);
   U18066 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_9_port, A2 => n11833, ZN 
                           => N95);
   U18067 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_10_port, A2 => n11834, ZN
                           => N96);
   U18068 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_11_port, A2 => n11834, ZN
                           => N97);
   U18069 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_12_port, A2 => n11835, ZN
                           => N98);
   U18070 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_13_port, A2 => n11836, ZN
                           => N99);
   U18071 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_14_port, A2 => n11667, ZN
                           => N100);
   U18072 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_15_port, A2 => n11667, ZN
                           => N101);
   U18073 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_16_port, A2 => n11668, ZN
                           => N102);
   U18074 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_17_port, A2 => n11669, ZN
                           => N103);
   U18075 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_18_port, A2 => n11670, ZN
                           => N104);
   U18076 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_19_port, A2 => n11671, ZN
                           => N105);
   U18077 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_20_port, A2 => n11672, ZN
                           => N106);
   U18078 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_21_port, A2 => n11673, ZN
                           => N107);
   U18079 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_22_port, A2 => n11674, ZN
                           => N108);
   U18080 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_23_port, A2 => n11675, ZN
                           => N109);
   U18081 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_24_port, A2 => n11676, ZN
                           => N110);
   U18082 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_25_port, A2 => n11677, ZN
                           => N111);
   U18083 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_26_port, A2 => n11678, ZN
                           => N112);
   U18084 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_27_port, A2 => n11678, ZN
                           => N113);
   U18085 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_28_port, A2 => n11679, ZN
                           => N114);
   U18086 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_29_port, A2 => n11680, ZN
                           => N115);
   U18087 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_30_port, A2 => n11681, ZN
                           => N116);
   U18088 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_31_port, A2 => n11682, ZN
                           => N117);
   U18089 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_32_port, A2 => n11683, ZN
                           => N118);
   U18090 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_33_port, A2 => n11684, ZN
                           => N119);
   U18091 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_34_port, A2 => n11685, ZN
                           => N120);
   U18092 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_35_port, A2 => n11686, ZN
                           => N121);
   U18093 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_36_port, A2 => n11687, ZN
                           => N122);
   U18094 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_37_port, A2 => n11688, ZN
                           => N123);
   U18095 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_38_port, A2 => n11689, ZN
                           => N124);
   U18096 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_39_port, A2 => n11689, ZN
                           => N125);
   U18097 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_40_port, A2 => n11690, ZN
                           => N126);
   U18098 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_41_port, A2 => n11691, ZN
                           => N127);
   U18099 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_42_port, A2 => n11692, ZN
                           => N128);
   U18100 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_43_port, A2 => n11693, ZN
                           => N129);
   U18101 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_44_port, A2 => n11694, ZN
                           => N130);
   U18102 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_45_port, A2 => n11695, ZN
                           => N131);
   U18103 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_46_port, A2 => n11696, ZN
                           => N132);
   U18104 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_47_port, A2 => n11697, ZN
                           => N133);
   U18105 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_48_port, A2 => n11698, ZN
                           => N134);
   U18106 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_49_port, A2 => n11699, ZN
                           => N135);
   U18107 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_50_port, A2 => n11700, ZN
                           => N136);
   U18108 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_51_port, A2 => n11700, ZN
                           => N137);
   U18109 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_52_port, A2 => n11701, ZN
                           => N138);
   U18110 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_53_port, A2 => n11702, ZN
                           => N139);
   U18111 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_54_port, A2 => n11703, ZN
                           => N140);
   U18112 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_55_port, A2 => n11704, ZN
                           => N141);
   U18113 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_56_port, A2 => n11705, ZN
                           => N142);
   U18114 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_57_port, A2 => n11706, ZN
                           => N143);
   U18115 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_58_port, A2 => n11707, ZN
                           => N144);
   U18116 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_59_port, A2 => n11708, ZN
                           => N145);
   U18117 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_60_port, A2 => n11709, ZN
                           => N146);
   U18118 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_61_port, A2 => n11710, ZN
                           => N147);
   U18119 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_62_port, A2 => n11711, ZN
                           => N148);
   U18120 : AND2_X1 port map( A1 => NEXT_REGISTERS_30_63_port, A2 => n11711, ZN
                           => N149);
   U18121 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_0_port, A2 => n11712, ZN 
                           => N150);
   U18122 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_1_port, A2 => n11713, ZN 
                           => N151);
   U18123 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_2_port, A2 => n11714, ZN 
                           => N152);
   U18124 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_3_port, A2 => n11715, ZN 
                           => N153);
   U18125 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_4_port, A2 => n11716, ZN 
                           => N154);
   U18126 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_5_port, A2 => n11717, ZN 
                           => N155);
   U18127 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_6_port, A2 => n11718, ZN 
                           => N156);
   U18128 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_7_port, A2 => n11719, ZN 
                           => N157);
   U18129 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_8_port, A2 => n11720, ZN 
                           => N158);
   U18130 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_9_port, A2 => n11721, ZN 
                           => N159);
   U18131 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_10_port, A2 => n11722, ZN
                           => N160);
   U18132 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_11_port, A2 => n11722, ZN
                           => N161);
   U18133 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_12_port, A2 => n11723, ZN
                           => N162);
   U18134 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_13_port, A2 => n11724, ZN
                           => N163);
   U18135 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_14_port, A2 => n11725, ZN
                           => N164);
   U18136 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_15_port, A2 => n11726, ZN
                           => N165);
   U18137 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_16_port, A2 => n11727, ZN
                           => N166);
   U18138 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_17_port, A2 => n11728, ZN
                           => N167);
   U18139 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_18_port, A2 => n11729, ZN
                           => N168);
   U18140 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_19_port, A2 => n11730, ZN
                           => N169);
   U18141 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_20_port, A2 => n11731, ZN
                           => N170);
   U18142 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_21_port, A2 => n11732, ZN
                           => N171);
   U18143 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_22_port, A2 => n11733, ZN
                           => N172);
   U18144 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_23_port, A2 => n11733, ZN
                           => N173);
   U18145 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_24_port, A2 => n11734, ZN
                           => N174);
   U18146 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_25_port, A2 => n11735, ZN
                           => N175);
   U18147 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_26_port, A2 => n11736, ZN
                           => N176);
   U18148 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_27_port, A2 => n11737, ZN
                           => N177);
   U18149 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_28_port, A2 => n11738, ZN
                           => N178);
   U18150 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_29_port, A2 => n11739, ZN
                           => N179);
   U18151 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_30_port, A2 => n11740, ZN
                           => N180);
   U18152 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_31_port, A2 => n11741, ZN
                           => N181);
   U18153 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_32_port, A2 => n11742, ZN
                           => N182);
   U18154 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_33_port, A2 => n11743, ZN
                           => N183);
   U18155 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_34_port, A2 => n11744, ZN
                           => N184);
   U18156 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_35_port, A2 => n11744, ZN
                           => N185);
   U18157 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_36_port, A2 => n11745, ZN
                           => N186);
   U18158 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_37_port, A2 => n11746, ZN
                           => N187);
   U18159 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_38_port, A2 => n11747, ZN
                           => N188);
   U18160 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_39_port, A2 => n11748, ZN
                           => N189);
   U18161 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_40_port, A2 => n11749, ZN
                           => N190);
   U18162 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_41_port, A2 => n11750, ZN
                           => N191);
   U18163 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_42_port, A2 => n11751, ZN
                           => N192);
   U18164 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_43_port, A2 => n11752, ZN
                           => N193);
   U18165 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_44_port, A2 => n11753, ZN
                           => N194);
   U18166 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_45_port, A2 => n11754, ZN
                           => N195);
   U18167 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_46_port, A2 => n11755, ZN
                           => N196);
   U18168 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_47_port, A2 => n11755, ZN
                           => N197);
   U18169 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_48_port, A2 => n11756, ZN
                           => N198);
   U18170 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_49_port, A2 => n11757, ZN
                           => N199);
   U18171 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_50_port, A2 => n11758, ZN
                           => N200);
   U18172 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_51_port, A2 => n11759, ZN
                           => N201);
   U18173 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_52_port, A2 => n11760, ZN
                           => N202);
   U18174 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_53_port, A2 => n11761, ZN
                           => N203);
   U18175 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_54_port, A2 => n11762, ZN
                           => N204);
   U18176 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_55_port, A2 => n11763, ZN
                           => N205);
   U18177 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_56_port, A2 => n11764, ZN
                           => N206);
   U18178 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_57_port, A2 => n11765, ZN
                           => N207);
   U18179 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_58_port, A2 => n11765, ZN
                           => N208);
   U18180 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_59_port, A2 => n11765, ZN
                           => N209);
   U18181 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_60_port, A2 => n11765, ZN
                           => N210);
   U18182 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_61_port, A2 => n11765, ZN
                           => N211);
   U18183 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_62_port, A2 => n11765, ZN
                           => N212);
   U18184 : AND2_X1 port map( A1 => NEXT_REGISTERS_29_63_port, A2 => n11765, ZN
                           => N213);
   U18185 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_0_port, A2 => n11765, ZN 
                           => N214);
   U18186 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_1_port, A2 => n11765, ZN 
                           => N215);
   U18187 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_2_port, A2 => n11765, ZN 
                           => N216);
   U18188 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_3_port, A2 => n11765, ZN 
                           => N217);
   U18189 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_4_port, A2 => n11766, ZN 
                           => N218);
   U18190 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_5_port, A2 => n11766, ZN 
                           => N219);
   U18191 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_6_port, A2 => n11766, ZN 
                           => N220);
   U18192 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_7_port, A2 => n11766, ZN 
                           => N221);
   U18193 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_8_port, A2 => n11766, ZN 
                           => N222);
   U18194 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_9_port, A2 => n11766, ZN 
                           => N223);
   U18195 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_10_port, A2 => n11766, ZN
                           => N224);
   U18196 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_11_port, A2 => n11766, ZN
                           => N225);
   U18197 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_12_port, A2 => n11766, ZN
                           => N226);
   U18198 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_13_port, A2 => n11766, ZN
                           => N227);
   U18199 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_14_port, A2 => n11766, ZN
                           => N228);
   U18200 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_15_port, A2 => n11767, ZN
                           => N229);
   U18201 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_16_port, A2 => n11767, ZN
                           => N230);
   U18202 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_17_port, A2 => n11767, ZN
                           => N231);
   U18203 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_18_port, A2 => n11767, ZN
                           => N232);
   U18204 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_19_port, A2 => n11767, ZN
                           => N233);
   U18205 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_20_port, A2 => n11767, ZN
                           => N234);
   U18206 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_21_port, A2 => n11767, ZN
                           => N235);
   U18207 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_22_port, A2 => n11767, ZN
                           => N236);
   U18208 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_23_port, A2 => n11767, ZN
                           => N237);
   U18209 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_24_port, A2 => n11767, ZN
                           => N238);
   U18210 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_25_port, A2 => n11767, ZN
                           => N239);
   U18211 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_26_port, A2 => n11768, ZN
                           => N240);
   U18212 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_27_port, A2 => n11768, ZN
                           => N241);
   U18213 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_28_port, A2 => n11768, ZN
                           => N242);
   U18214 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_29_port, A2 => n11768, ZN
                           => N243);
   U18215 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_30_port, A2 => n11768, ZN
                           => N244);
   U18216 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_31_port, A2 => n11768, ZN
                           => N245);
   U18217 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_32_port, A2 => n11768, ZN
                           => N246);
   U18218 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_33_port, A2 => n11768, ZN
                           => N247);
   U18219 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_34_port, A2 => n11768, ZN
                           => N248);
   U18220 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_35_port, A2 => n11768, ZN
                           => N249);
   U18221 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_36_port, A2 => n11769, ZN
                           => N250);
   U18222 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_37_port, A2 => n11769, ZN
                           => N251);
   U18223 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_38_port, A2 => n11769, ZN
                           => N252);
   U18224 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_39_port, A2 => n11769, ZN
                           => N253);
   U18225 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_40_port, A2 => n11769, ZN
                           => N254);
   U18226 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_41_port, A2 => n11769, ZN
                           => N255);
   U18227 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_42_port, A2 => n11769, ZN
                           => N256);
   U18228 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_43_port, A2 => n11769, ZN
                           => N257);
   U18229 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_44_port, A2 => n11769, ZN
                           => N258);
   U18230 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_45_port, A2 => n11769, ZN
                           => N259);
   U18231 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_46_port, A2 => n11769, ZN
                           => N260);
   U18232 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_47_port, A2 => n11770, ZN
                           => N261);
   U18233 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_48_port, A2 => n11770, ZN
                           => N262);
   U18234 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_49_port, A2 => n11770, ZN
                           => N263);
   U18235 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_50_port, A2 => n11770, ZN
                           => N264);
   U18236 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_51_port, A2 => n11770, ZN
                           => N265);
   U18237 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_52_port, A2 => n11770, ZN
                           => N266);
   U18238 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_53_port, A2 => n11770, ZN
                           => N267);
   U18239 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_54_port, A2 => n11770, ZN
                           => N268);
   U18240 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_55_port, A2 => n11770, ZN
                           => N269);
   U18241 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_56_port, A2 => n11770, ZN
                           => N270);
   U18242 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_57_port, A2 => n11770, ZN
                           => N271);
   U18243 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_58_port, A2 => n11771, ZN
                           => N272);
   U18244 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_59_port, A2 => n11771, ZN
                           => N273);
   U18245 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_60_port, A2 => n11771, ZN
                           => N274);
   U18246 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_61_port, A2 => n11771, ZN
                           => N275);
   U18247 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_62_port, A2 => n11771, ZN
                           => N276);
   U18248 : AND2_X1 port map( A1 => NEXT_REGISTERS_28_63_port, A2 => n11771, ZN
                           => N277);
   U18249 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_0_port, A2 => n11771, ZN 
                           => N278);
   U18250 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_1_port, A2 => n11771, ZN 
                           => N279);
   U18251 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_2_port, A2 => n11771, ZN 
                           => N280);
   U18252 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_3_port, A2 => n11771, ZN 
                           => N281);
   U18253 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_4_port, A2 => n11771, ZN 
                           => N282);
   U18254 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_5_port, A2 => n11772, ZN 
                           => N283);
   U18255 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_6_port, A2 => n11772, ZN 
                           => N284);
   U18256 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_7_port, A2 => n11772, ZN 
                           => N285);
   U18257 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_8_port, A2 => n11772, ZN 
                           => N286);
   U18258 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_9_port, A2 => n11772, ZN 
                           => N287);
   U18259 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_10_port, A2 => n11772, ZN
                           => N288);
   U18260 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_11_port, A2 => n11772, ZN
                           => N289);
   U18261 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_12_port, A2 => n11772, ZN
                           => N290);
   U18262 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_13_port, A2 => n11772, ZN
                           => N291);
   U18263 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_14_port, A2 => n11772, ZN
                           => N292);
   U18264 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_15_port, A2 => n11772, ZN
                           => N293);
   U18265 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_16_port, A2 => n11773, ZN
                           => N294);
   U18266 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_17_port, A2 => n11773, ZN
                           => N295);
   U18267 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_18_port, A2 => n11773, ZN
                           => N296);
   U18268 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_19_port, A2 => n11773, ZN
                           => N297);
   U18269 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_20_port, A2 => n11773, ZN
                           => N298);
   U18270 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_21_port, A2 => n11773, ZN
                           => N299);
   U18271 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_22_port, A2 => n11773, ZN
                           => N300);
   U18272 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_23_port, A2 => n11773, ZN
                           => N301);
   U18273 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_24_port, A2 => n11773, ZN
                           => N302);
   U18274 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_25_port, A2 => n11773, ZN
                           => N303);
   U18275 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_26_port, A2 => n11773, ZN
                           => N304);
   U18276 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_27_port, A2 => n11774, ZN
                           => N305);
   U18277 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_28_port, A2 => n11774, ZN
                           => N306);
   U18278 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_29_port, A2 => n11774, ZN
                           => N307);
   U18279 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_30_port, A2 => n11774, ZN
                           => N308);
   U18280 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_31_port, A2 => n11774, ZN
                           => N309);
   U18281 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_32_port, A2 => n11774, ZN
                           => N310);
   U18282 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_33_port, A2 => n11774, ZN
                           => N311);
   U18283 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_34_port, A2 => n11774, ZN
                           => N312);
   U18284 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_35_port, A2 => n11774, ZN
                           => N313);
   U18285 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_36_port, A2 => n11774, ZN
                           => N314);
   U18286 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_37_port, A2 => n11774, ZN
                           => N315);
   U18287 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_38_port, A2 => n11775, ZN
                           => N316);
   U18288 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_39_port, A2 => n11775, ZN
                           => N317);
   U18289 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_40_port, A2 => n11775, ZN
                           => N318);
   U18290 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_41_port, A2 => n11775, ZN
                           => N319);
   U18291 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_42_port, A2 => n11775, ZN
                           => N320);
   U18292 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_43_port, A2 => n11775, ZN
                           => N321);
   U18293 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_44_port, A2 => n11775, ZN
                           => N322);
   U18294 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_45_port, A2 => n11775, ZN
                           => N323);
   U18295 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_46_port, A2 => n11775, ZN
                           => N324);
   U18296 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_47_port, A2 => n11775, ZN
                           => N325);
   U18297 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_48_port, A2 => n11775, ZN
                           => N326);
   U18298 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_49_port, A2 => n11776, ZN
                           => N327);
   U18299 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_50_port, A2 => n11776, ZN
                           => N328);
   U18300 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_51_port, A2 => n11776, ZN
                           => N329);
   U18301 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_52_port, A2 => n11776, ZN
                           => N330);
   U18302 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_53_port, A2 => n11776, ZN
                           => N331);
   U18303 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_54_port, A2 => n11776, ZN
                           => N332);
   U18304 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_55_port, A2 => n11776, ZN
                           => N333);
   U18305 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_56_port, A2 => n11776, ZN
                           => N334);
   U18306 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_57_port, A2 => n11776, ZN
                           => N335);
   U18307 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_58_port, A2 => n11776, ZN
                           => N336);
   U18308 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_59_port, A2 => n11776, ZN
                           => N337);
   U18309 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_60_port, A2 => n11777, ZN
                           => N338);
   U18310 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_61_port, A2 => n11777, ZN
                           => N339);
   U18311 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_62_port, A2 => n11777, ZN
                           => N340);
   U18312 : AND2_X1 port map( A1 => NEXT_REGISTERS_27_63_port, A2 => n11777, ZN
                           => N341);
   U18313 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_0_port, A2 => n11777, ZN 
                           => N342);
   U18314 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_1_port, A2 => n11777, ZN 
                           => N343);
   U18315 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_2_port, A2 => n11777, ZN 
                           => N344);
   U18316 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_3_port, A2 => n11777, ZN 
                           => N345);
   U18317 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_4_port, A2 => n11777, ZN 
                           => N346);
   U18318 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_5_port, A2 => n11777, ZN 
                           => N347);
   U18319 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_6_port, A2 => n11777, ZN 
                           => N348);
   U18320 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_7_port, A2 => n11778, ZN 
                           => N349);
   U18321 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_8_port, A2 => n11778, ZN 
                           => N350);
   U18322 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_9_port, A2 => n11778, ZN 
                           => N351);
   U18323 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_10_port, A2 => n11778, ZN
                           => N352);
   U18324 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_11_port, A2 => n11778, ZN
                           => N353);
   U18325 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_12_port, A2 => n11778, ZN
                           => N354);
   U18326 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_13_port, A2 => n11778, ZN
                           => N355);
   U18327 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_14_port, A2 => n11778, ZN
                           => N356);
   U18328 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_15_port, A2 => n11778, ZN
                           => N357);
   U18329 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_16_port, A2 => n11778, ZN
                           => N358);
   U18330 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_17_port, A2 => n11778, ZN
                           => N359);
   U18331 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_18_port, A2 => n11779, ZN
                           => N360);
   U18332 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_19_port, A2 => n11779, ZN
                           => N361);
   U18333 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_20_port, A2 => n11779, ZN
                           => N362);
   U18334 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_21_port, A2 => n11779, ZN
                           => N363);
   U18335 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_22_port, A2 => n11779, ZN
                           => N364);
   U18336 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_23_port, A2 => n11779, ZN
                           => N365);
   U18337 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_24_port, A2 => n11779, ZN
                           => N366);
   U18338 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_25_port, A2 => n11779, ZN
                           => N367);
   U18339 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_26_port, A2 => n11779, ZN
                           => N368);
   U18340 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_27_port, A2 => n11779, ZN
                           => N369);
   U18341 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_28_port, A2 => n11780, ZN
                           => N370);
   U18342 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_29_port, A2 => n11780, ZN
                           => N371);
   U18343 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_30_port, A2 => n11780, ZN
                           => N372);
   U18344 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_31_port, A2 => n11780, ZN
                           => N373);
   U18345 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_32_port, A2 => n11780, ZN
                           => N374);
   U18346 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_33_port, A2 => n11780, ZN
                           => N375);
   U18347 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_34_port, A2 => n11780, ZN
                           => N376);
   U18348 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_35_port, A2 => n11780, ZN
                           => N377);
   U18349 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_36_port, A2 => n11780, ZN
                           => N378);
   U18350 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_37_port, A2 => n11780, ZN
                           => N379);
   U18351 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_38_port, A2 => n11780, ZN
                           => N380);
   U18352 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_39_port, A2 => n11781, ZN
                           => N381);
   U18353 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_40_port, A2 => n11781, ZN
                           => N382);
   U18354 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_41_port, A2 => n11781, ZN
                           => N383);
   U18355 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_42_port, A2 => n11781, ZN
                           => N384);
   U18356 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_43_port, A2 => n11781, ZN
                           => N385);
   U18357 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_44_port, A2 => n11781, ZN
                           => N386);
   U18358 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_45_port, A2 => n11781, ZN
                           => N387);
   U18359 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_46_port, A2 => n11781, ZN
                           => N388);
   U18360 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_47_port, A2 => n11781, ZN
                           => N389);
   U18361 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_48_port, A2 => n11781, ZN
                           => N390);
   U18362 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_49_port, A2 => n11781, ZN
                           => N391);
   U18363 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_50_port, A2 => n11782, ZN
                           => N392);
   U18364 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_51_port, A2 => n11782, ZN
                           => N393);
   U18365 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_52_port, A2 => n11782, ZN
                           => N394);
   U18366 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_53_port, A2 => n11782, ZN
                           => N395);
   U18367 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_54_port, A2 => n11782, ZN
                           => N396);
   U18368 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_55_port, A2 => n11782, ZN
                           => N397);
   U18369 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_56_port, A2 => n11782, ZN
                           => N398);
   U18370 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_57_port, A2 => n11782, ZN
                           => N399);
   U18371 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_58_port, A2 => n11782, ZN
                           => N400);
   U18372 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_59_port, A2 => n11782, ZN
                           => N401);
   U18373 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_60_port, A2 => n11782, ZN
                           => N402);
   U18374 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_61_port, A2 => n11783, ZN
                           => N403);
   U18375 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_62_port, A2 => n11783, ZN
                           => N404);
   U18376 : AND2_X1 port map( A1 => NEXT_REGISTERS_26_63_port, A2 => n11783, ZN
                           => N405);
   U18377 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_0_port, A2 => n11783, ZN 
                           => N406);
   U18378 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_1_port, A2 => n11783, ZN 
                           => N407);
   U18379 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_2_port, A2 => n11783, ZN 
                           => N408);
   U18380 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_3_port, A2 => n11783, ZN 
                           => N409);
   U18381 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_4_port, A2 => n11783, ZN 
                           => N410);
   U18382 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_5_port, A2 => n11783, ZN 
                           => N411);
   U18383 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_6_port, A2 => n11783, ZN 
                           => N412);
   U18384 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_7_port, A2 => n11783, ZN 
                           => N413);
   U18385 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_8_port, A2 => n11784, ZN 
                           => N414);
   U18386 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_9_port, A2 => n11784, ZN 
                           => N415);
   U18387 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_10_port, A2 => n11784, ZN
                           => N416);
   U18388 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_11_port, A2 => n11784, ZN
                           => N417);
   U18389 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_12_port, A2 => n11784, ZN
                           => N418);
   U18390 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_13_port, A2 => n11784, ZN
                           => N419);
   U18391 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_14_port, A2 => n11784, ZN
                           => N420);
   U18392 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_15_port, A2 => n11784, ZN
                           => N421);
   U18393 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_16_port, A2 => n11784, ZN
                           => N422);
   U18394 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_17_port, A2 => n11784, ZN
                           => N423);
   U18395 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_18_port, A2 => n11784, ZN
                           => N424);
   U18396 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_19_port, A2 => n11785, ZN
                           => N425);
   U18397 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_20_port, A2 => n11785, ZN
                           => N426);
   U18398 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_21_port, A2 => n11785, ZN
                           => N427);
   U18399 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_22_port, A2 => n11785, ZN
                           => N428);
   U18400 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_23_port, A2 => n11785, ZN
                           => N429);
   U18401 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_24_port, A2 => n11785, ZN
                           => N430);
   U18402 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_25_port, A2 => n11785, ZN
                           => N431);
   U18403 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_26_port, A2 => n11785, ZN
                           => N432);
   U18404 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_27_port, A2 => n11785, ZN
                           => N433);
   U18405 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_28_port, A2 => n11785, ZN
                           => N434);
   U18406 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_29_port, A2 => n11785, ZN
                           => N435);
   U18407 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_30_port, A2 => n11786, ZN
                           => N436);
   U18408 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_31_port, A2 => n11786, ZN
                           => N437);
   U18409 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_32_port, A2 => n11786, ZN
                           => N438);
   U18410 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_33_port, A2 => n11786, ZN
                           => N439);
   U18411 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_34_port, A2 => n11786, ZN
                           => N440);
   U18412 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_35_port, A2 => n11786, ZN
                           => N441);
   U18413 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_36_port, A2 => n11786, ZN
                           => N442);
   U18414 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_37_port, A2 => n11786, ZN
                           => N443);
   U18415 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_38_port, A2 => n11786, ZN
                           => N444);
   U18416 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_39_port, A2 => n11786, ZN
                           => N445);
   U18417 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_40_port, A2 => n11786, ZN
                           => N446);
   U18418 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_41_port, A2 => n11787, ZN
                           => N447);
   U18419 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_42_port, A2 => n11787, ZN
                           => N448);
   U18420 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_43_port, A2 => n11787, ZN
                           => N449);
   U18421 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_44_port, A2 => n11787, ZN
                           => N450);
   U18422 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_45_port, A2 => n11787, ZN
                           => N451);
   U18423 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_46_port, A2 => n11787, ZN
                           => N452);
   U18424 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_47_port, A2 => n11787, ZN
                           => N453);
   U18425 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_48_port, A2 => n11787, ZN
                           => N454);
   U18426 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_49_port, A2 => n11787, ZN
                           => N455);
   U18427 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_50_port, A2 => n11787, ZN
                           => N456);
   U18428 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_51_port, A2 => n11787, ZN
                           => N457);
   U18429 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_52_port, A2 => n11788, ZN
                           => N458);
   U18430 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_53_port, A2 => n11788, ZN
                           => N459);
   U18431 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_54_port, A2 => n11788, ZN
                           => N460);
   U18432 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_55_port, A2 => n11788, ZN
                           => N461);
   U18433 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_56_port, A2 => n11788, ZN
                           => N462);
   U18434 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_57_port, A2 => n11788, ZN
                           => N463);
   U18435 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_58_port, A2 => n11788, ZN
                           => N464);
   U18436 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_59_port, A2 => n11788, ZN
                           => N465);
   U18437 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_60_port, A2 => n11788, ZN
                           => N466);
   U18438 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_61_port, A2 => n11788, ZN
                           => N467);
   U18439 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_62_port, A2 => n11788, ZN
                           => N468);
   U18440 : AND2_X1 port map( A1 => NEXT_REGISTERS_25_63_port, A2 => n11789, ZN
                           => N469);
   U18441 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_0_port, A2 => n11789, ZN 
                           => N470);
   U18442 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_1_port, A2 => n11789, ZN 
                           => N471);
   U18443 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_2_port, A2 => n11789, ZN 
                           => N472);
   U18444 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_3_port, A2 => n11789, ZN 
                           => N473);
   U18445 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_4_port, A2 => n11789, ZN 
                           => N474);
   U18446 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_5_port, A2 => n11789, ZN 
                           => N475);
   U18447 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_6_port, A2 => n11789, ZN 
                           => N476);
   U18448 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_7_port, A2 => n11789, ZN 
                           => N477);
   U18449 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_8_port, A2 => n11789, ZN 
                           => N478);
   U18450 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_9_port, A2 => n11789, ZN 
                           => N479);
   U18451 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_10_port, A2 => n11790, ZN
                           => N480);
   U18452 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_11_port, A2 => n11790, ZN
                           => N481);
   U18453 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_12_port, A2 => n11790, ZN
                           => N482);
   U18454 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_13_port, A2 => n11790, ZN
                           => N483);
   U18455 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_14_port, A2 => n11790, ZN
                           => N484);
   U18456 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_15_port, A2 => n11790, ZN
                           => N485);
   U18457 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_16_port, A2 => n11790, ZN
                           => N486);
   U18458 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_17_port, A2 => n11790, ZN
                           => N487);
   U18459 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_18_port, A2 => n11790, ZN
                           => N488);
   U18460 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_19_port, A2 => n11790, ZN
                           => N489);
   U18461 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_20_port, A2 => n11791, ZN
                           => N490);
   U18462 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_21_port, A2 => n11791, ZN
                           => N491);
   U18463 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_22_port, A2 => n11791, ZN
                           => N492);
   U18464 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_23_port, A2 => n11791, ZN
                           => N493);
   U18465 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_24_port, A2 => n11791, ZN
                           => N494);
   U18466 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_25_port, A2 => n11791, ZN
                           => N495);
   U18467 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_26_port, A2 => n11791, ZN
                           => N496);
   U18468 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_27_port, A2 => n11791, ZN
                           => N497);
   U18469 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_28_port, A2 => n11791, ZN
                           => N498);
   U18470 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_29_port, A2 => n11791, ZN
                           => N499);
   U18471 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_30_port, A2 => n11791, ZN
                           => N500);
   U18472 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_31_port, A2 => n11792, ZN
                           => N501);
   U18473 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_32_port, A2 => n11792, ZN
                           => N502);
   U18474 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_33_port, A2 => n11792, ZN
                           => N503);
   U18475 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_34_port, A2 => n11792, ZN
                           => N504);
   U18476 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_35_port, A2 => n11792, ZN
                           => N505);
   U18477 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_36_port, A2 => n11792, ZN
                           => N506);
   U18478 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_37_port, A2 => n11792, ZN
                           => N507);
   U18479 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_38_port, A2 => n11792, ZN
                           => N508);
   U18480 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_39_port, A2 => n11792, ZN
                           => N509);
   U18481 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_40_port, A2 => n11792, ZN
                           => N510);
   U18482 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_41_port, A2 => n11792, ZN
                           => N511);
   U18483 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_42_port, A2 => n11793, ZN
                           => N512);
   U18484 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_43_port, A2 => n11793, ZN
                           => N513);
   U18485 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_44_port, A2 => n11793, ZN
                           => N514);
   U18486 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_45_port, A2 => n11793, ZN
                           => N515);
   U18487 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_46_port, A2 => n11793, ZN
                           => N516);
   U18488 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_47_port, A2 => n11793, ZN
                           => N517);
   U18489 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_48_port, A2 => n11793, ZN
                           => N518);
   U18490 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_49_port, A2 => n11793, ZN
                           => N519);
   U18491 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_50_port, A2 => n11793, ZN
                           => N520);
   U18492 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_51_port, A2 => n11793, ZN
                           => N521);
   U18493 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_52_port, A2 => n11793, ZN
                           => N522);
   U18494 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_53_port, A2 => n11794, ZN
                           => N523);
   U18495 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_54_port, A2 => n11794, ZN
                           => N524);
   U18496 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_55_port, A2 => n11794, ZN
                           => N525);
   U18497 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_56_port, A2 => n11794, ZN
                           => N526);
   U18498 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_57_port, A2 => n11794, ZN
                           => N527);
   U18499 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_58_port, A2 => n11794, ZN
                           => N528);
   U18500 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_59_port, A2 => n11794, ZN
                           => N529);
   U18501 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_60_port, A2 => n11794, ZN
                           => N530);
   U18502 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_61_port, A2 => n11794, ZN
                           => N531);
   U18503 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_62_port, A2 => n11794, ZN
                           => N532);
   U18504 : AND2_X1 port map( A1 => NEXT_REGISTERS_24_63_port, A2 => n11794, ZN
                           => N533);
   U18505 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_0_port, A2 => n11795, ZN 
                           => N534);
   U18506 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_1_port, A2 => n11795, ZN 
                           => N535);
   U18507 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_2_port, A2 => n11795, ZN 
                           => N536);
   U18508 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_3_port, A2 => n11795, ZN 
                           => N537);
   U18509 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_4_port, A2 => n11795, ZN 
                           => N538);
   U18510 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_5_port, A2 => n11795, ZN 
                           => N539);
   U18511 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_6_port, A2 => n11795, ZN 
                           => N540);
   U18512 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_7_port, A2 => n11795, ZN 
                           => N541);
   U18513 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_8_port, A2 => n11795, ZN 
                           => N542);
   U18514 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_9_port, A2 => n11795, ZN 
                           => N543);
   U18515 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_10_port, A2 => n11795, ZN
                           => N544);
   U18516 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_11_port, A2 => n11796, ZN
                           => N545);
   U18517 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_12_port, A2 => n11796, ZN
                           => N546);
   U18518 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_13_port, A2 => n11796, ZN
                           => N547);
   U18519 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_14_port, A2 => n11796, ZN
                           => N548);
   U18520 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_15_port, A2 => n11796, ZN
                           => N549);
   U18521 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_16_port, A2 => n11796, ZN
                           => N550);
   U18522 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_17_port, A2 => n11796, ZN
                           => N551);
   U18523 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_18_port, A2 => n11796, ZN
                           => N552);
   U18524 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_19_port, A2 => n11796, ZN
                           => N553);
   U18525 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_20_port, A2 => n11796, ZN
                           => N554);
   U18526 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_21_port, A2 => n11796, ZN
                           => N555);
   U18527 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_22_port, A2 => n11797, ZN
                           => N556);
   U18528 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_23_port, A2 => n11797, ZN
                           => N557);
   U18529 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_24_port, A2 => n11797, ZN
                           => N558);
   U18530 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_25_port, A2 => n11797, ZN
                           => N559);
   U18531 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_26_port, A2 => n11797, ZN
                           => N560);
   U18532 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_27_port, A2 => n11797, ZN
                           => N561);
   U18533 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_28_port, A2 => n11797, ZN
                           => N562);
   U18534 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_29_port, A2 => n11797, ZN
                           => N563);
   U18535 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_30_port, A2 => n11797, ZN
                           => N564);
   U18536 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_31_port, A2 => n11797, ZN
                           => N565);
   U18537 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_32_port, A2 => n11797, ZN
                           => N566);
   U18538 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_33_port, A2 => n11798, ZN
                           => N567);
   U18539 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_34_port, A2 => n11798, ZN
                           => N568);
   U18540 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_35_port, A2 => n11798, ZN
                           => N569);
   U18541 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_36_port, A2 => n11798, ZN
                           => N570);
   U18542 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_37_port, A2 => n11798, ZN
                           => N571);
   U18543 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_38_port, A2 => n11798, ZN
                           => N572);
   U18544 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_39_port, A2 => n11798, ZN
                           => N573);
   U18545 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_40_port, A2 => n11798, ZN
                           => N574);
   U18546 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_41_port, A2 => n11798, ZN
                           => N575);
   U18547 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_42_port, A2 => n11798, ZN
                           => N576);
   U18548 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_43_port, A2 => n11798, ZN
                           => N577);
   U18549 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_44_port, A2 => n11799, ZN
                           => N578);
   U18550 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_45_port, A2 => n11799, ZN
                           => N579);
   U18551 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_46_port, A2 => n11799, ZN
                           => N580);
   U18552 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_47_port, A2 => n11799, ZN
                           => N581);
   U18553 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_48_port, A2 => n11799, ZN
                           => N582);
   U18554 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_49_port, A2 => n11799, ZN
                           => N583);
   U18555 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_50_port, A2 => n11799, ZN
                           => N584);
   U18556 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_51_port, A2 => n11799, ZN
                           => N585);
   U18557 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_52_port, A2 => n11799, ZN
                           => N586);
   U18558 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_53_port, A2 => n11799, ZN
                           => N587);
   U18559 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_54_port, A2 => n11799, ZN
                           => N588);
   U18560 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_55_port, A2 => n11800, ZN
                           => N589);
   U18561 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_56_port, A2 => n11800, ZN
                           => N590);
   U18562 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_57_port, A2 => n11800, ZN
                           => N591);
   U18563 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_58_port, A2 => n11800, ZN
                           => N592);
   U18564 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_59_port, A2 => n11800, ZN
                           => N593);
   U18565 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_60_port, A2 => n11800, ZN
                           => N594);
   U18566 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_61_port, A2 => n11800, ZN
                           => N595);
   U18567 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_62_port, A2 => n11800, ZN
                           => N596);
   U18568 : AND2_X1 port map( A1 => NEXT_REGISTERS_23_63_port, A2 => n11800, ZN
                           => N597);
   U18569 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_0_port, A2 => n11800, ZN 
                           => N598);
   U18570 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_1_port, A2 => n11800, ZN 
                           => N599);
   U18571 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_2_port, A2 => n11801, ZN 
                           => N600);
   U18572 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_3_port, A2 => n11801, ZN 
                           => N601);
   U18573 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_4_port, A2 => n11801, ZN 
                           => N602);
   U18574 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_5_port, A2 => n11801, ZN 
                           => N603);
   U18575 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_6_port, A2 => n11801, ZN 
                           => N604);
   U18576 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_7_port, A2 => n11801, ZN 
                           => N605);
   U18577 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_8_port, A2 => n11801, ZN 
                           => N606);
   U18578 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_9_port, A2 => n11801, ZN 
                           => N607);
   U18579 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_10_port, A2 => n11801, ZN
                           => N608);
   U18580 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_11_port, A2 => n11801, ZN
                           => N609);
   U18581 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_12_port, A2 => n11802, ZN
                           => N610);
   U18582 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_13_port, A2 => n11802, ZN
                           => N611);
   U18583 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_14_port, A2 => n11802, ZN
                           => N612);
   U18584 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_15_port, A2 => n11802, ZN
                           => N613);
   U18585 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_16_port, A2 => n11802, ZN
                           => N614);
   U18586 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_17_port, A2 => n11802, ZN
                           => N615);
   U18587 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_18_port, A2 => n11802, ZN
                           => N616);
   U18588 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_19_port, A2 => n11802, ZN
                           => N617);
   U18589 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_20_port, A2 => n11802, ZN
                           => N618);
   U18590 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_21_port, A2 => n11802, ZN
                           => N619);
   U18591 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_22_port, A2 => n11802, ZN
                           => N620);
   U18592 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_23_port, A2 => n11803, ZN
                           => N621);
   U18593 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_24_port, A2 => n11803, ZN
                           => N622);
   U18594 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_25_port, A2 => n11803, ZN
                           => N623);
   U18595 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_26_port, A2 => n11803, ZN
                           => N624);
   U18596 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_27_port, A2 => n11803, ZN
                           => N625);
   U18597 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_28_port, A2 => n11803, ZN
                           => N626);
   U18598 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_29_port, A2 => n11803, ZN
                           => N627);
   U18599 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_30_port, A2 => n11803, ZN
                           => N628);
   U18600 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_31_port, A2 => n11803, ZN
                           => N629);
   U18601 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_32_port, A2 => n11803, ZN
                           => N630);
   U18602 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_33_port, A2 => n11803, ZN
                           => N631);
   U18603 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_34_port, A2 => n11804, ZN
                           => N632);
   U18604 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_35_port, A2 => n11804, ZN
                           => N633);
   U18605 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_36_port, A2 => n11804, ZN
                           => N634);
   U18606 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_37_port, A2 => n11804, ZN
                           => N635);
   U18607 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_38_port, A2 => n11804, ZN
                           => N636);
   U18608 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_39_port, A2 => n11804, ZN
                           => N637);
   U18609 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_40_port, A2 => n11804, ZN
                           => N638);
   U18610 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_41_port, A2 => n11804, ZN
                           => N639);
   U18611 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_42_port, A2 => n11804, ZN
                           => N640);
   U18612 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_43_port, A2 => n11804, ZN
                           => N641);
   U18613 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_44_port, A2 => n11804, ZN
                           => N642);
   U18614 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_45_port, A2 => n11805, ZN
                           => N643);
   U18615 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_46_port, A2 => n11805, ZN
                           => N644);
   U18616 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_47_port, A2 => n11805, ZN
                           => N645);
   U18617 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_48_port, A2 => n11805, ZN
                           => N646);
   U18618 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_49_port, A2 => n11805, ZN
                           => N647);
   U18619 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_50_port, A2 => n11805, ZN
                           => N648);
   U18620 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_51_port, A2 => n11805, ZN
                           => N649);
   U18621 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_52_port, A2 => n11805, ZN
                           => N650);
   U18622 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_53_port, A2 => n11805, ZN
                           => N651);
   U18623 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_54_port, A2 => n11805, ZN
                           => N652);
   U18624 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_55_port, A2 => n11805, ZN
                           => N653);
   U18625 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_56_port, A2 => n11806, ZN
                           => N654);
   U18626 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_57_port, A2 => n11806, ZN
                           => N655);
   U18627 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_58_port, A2 => n11806, ZN
                           => N656);
   U18628 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_59_port, A2 => n11806, ZN
                           => N657);
   U18629 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_60_port, A2 => n11806, ZN
                           => N658);
   U18630 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_61_port, A2 => n11806, ZN
                           => N659);
   U18631 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_62_port, A2 => n11806, ZN
                           => N660);
   U18632 : AND2_X1 port map( A1 => NEXT_REGISTERS_22_63_port, A2 => n11806, ZN
                           => N661);
   U18633 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_0_port, A2 => n11806, ZN 
                           => N662);
   U18634 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_1_port, A2 => n11806, ZN 
                           => N663);
   U18635 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_2_port, A2 => n11806, ZN 
                           => N664);
   U18636 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_3_port, A2 => n11807, ZN 
                           => N665);
   U18637 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_4_port, A2 => n11807, ZN 
                           => N666);
   U18638 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_5_port, A2 => n11807, ZN 
                           => N667);
   U18639 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_6_port, A2 => n11807, ZN 
                           => N668);
   U18640 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_7_port, A2 => n11807, ZN 
                           => N669);
   U18641 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_8_port, A2 => n11807, ZN 
                           => N670);
   U18642 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_9_port, A2 => n11807, ZN 
                           => N671);
   U18643 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_10_port, A2 => n11807, ZN
                           => N672);
   U18644 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_11_port, A2 => n11807, ZN
                           => N673);
   U18645 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_12_port, A2 => n11807, ZN
                           => N674);
   U18646 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_13_port, A2 => n11807, ZN
                           => N675);
   U18647 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_14_port, A2 => n11808, ZN
                           => N676);
   U18648 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_15_port, A2 => n11808, ZN
                           => N677);
   U18649 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_16_port, A2 => n11808, ZN
                           => N678);
   U18650 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_17_port, A2 => n11808, ZN
                           => N679);
   U18651 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_18_port, A2 => n11808, ZN
                           => N680);
   U18652 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_19_port, A2 => n11808, ZN
                           => N681);
   U18653 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_20_port, A2 => n11808, ZN
                           => N682);
   U18654 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_21_port, A2 => n11808, ZN
                           => N683);
   U18655 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_22_port, A2 => n11808, ZN
                           => N684);
   U18656 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_23_port, A2 => n11808, ZN
                           => N685);
   U18657 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_24_port, A2 => n11808, ZN
                           => N686);
   U18658 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_25_port, A2 => n11809, ZN
                           => N687);
   U18659 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_26_port, A2 => n11809, ZN
                           => N688);
   U18660 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_27_port, A2 => n11809, ZN
                           => N689);
   U18661 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_28_port, A2 => n11809, ZN
                           => N690);
   U18662 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_29_port, A2 => n11809, ZN
                           => N691);
   U18663 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_30_port, A2 => n11809, ZN
                           => N692);
   U18664 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_31_port, A2 => n11809, ZN
                           => N693);
   U18665 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_32_port, A2 => n11809, ZN
                           => N694);
   U18666 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_33_port, A2 => n11809, ZN
                           => N695);
   U18667 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_34_port, A2 => n11809, ZN
                           => N696);
   U18668 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_35_port, A2 => n11809, ZN
                           => N697);
   U18669 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_36_port, A2 => n11810, ZN
                           => N698);
   U18670 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_37_port, A2 => n11810, ZN
                           => N699);
   U18671 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_38_port, A2 => n11810, ZN
                           => N700);
   U18672 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_39_port, A2 => n11810, ZN
                           => N701);
   U18673 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_40_port, A2 => n11810, ZN
                           => N702);
   U18674 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_41_port, A2 => n11810, ZN
                           => N703);
   U18675 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_42_port, A2 => n11810, ZN
                           => N704);
   U18676 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_43_port, A2 => n11810, ZN
                           => N705);
   U18677 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_44_port, A2 => n11810, ZN
                           => N706);
   U18678 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_45_port, A2 => n11810, ZN
                           => N707);
   U18679 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_46_port, A2 => n11810, ZN
                           => N708);
   U18680 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_47_port, A2 => n11811, ZN
                           => N709);
   U18681 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_48_port, A2 => n11811, ZN
                           => N710);
   U18682 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_49_port, A2 => n11811, ZN
                           => N711);
   U18683 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_50_port, A2 => n11811, ZN
                           => N712);
   U18684 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_51_port, A2 => n11811, ZN
                           => N713);
   U18685 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_52_port, A2 => n11811, ZN
                           => N714);
   U18686 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_53_port, A2 => n11811, ZN
                           => N715);
   U18687 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_54_port, A2 => n11811, ZN
                           => N716);
   U18688 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_55_port, A2 => n11811, ZN
                           => N717);
   U18689 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_56_port, A2 => n11811, ZN
                           => N718);
   U18690 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_57_port, A2 => n11811, ZN
                           => N719);
   U18691 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_58_port, A2 => n11812, ZN
                           => N720);
   U18692 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_59_port, A2 => n11812, ZN
                           => N721);
   U18693 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_60_port, A2 => n11812, ZN
                           => N722);
   U18694 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_61_port, A2 => n11812, ZN
                           => N723);
   U18695 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_62_port, A2 => n11812, ZN
                           => N724);
   U18696 : AND2_X1 port map( A1 => NEXT_REGISTERS_21_63_port, A2 => n11812, ZN
                           => N725);
   U18697 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_0_port, A2 => n11812, ZN 
                           => N726);
   U18698 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_1_port, A2 => n11812, ZN 
                           => N727);
   U18699 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_2_port, A2 => n11812, ZN 
                           => N728);
   U18700 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_3_port, A2 => n11812, ZN 
                           => N729);
   U18701 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_4_port, A2 => n11813, ZN 
                           => N730);
   U18702 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_5_port, A2 => n11813, ZN 
                           => N731);
   U18703 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_6_port, A2 => n11813, ZN 
                           => N732);
   U18704 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_7_port, A2 => n11813, ZN 
                           => N733);
   U18705 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_8_port, A2 => n11813, ZN 
                           => N734);
   U18706 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_9_port, A2 => n11813, ZN 
                           => N735);
   U18707 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_10_port, A2 => n11813, ZN
                           => N736);
   U18708 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_11_port, A2 => n11813, ZN
                           => N737);
   U18709 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_12_port, A2 => n11813, ZN
                           => N738);
   U18710 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_13_port, A2 => n11813, ZN
                           => N739);
   U18711 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_14_port, A2 => n11813, ZN
                           => N740);
   U18712 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_15_port, A2 => n11814, ZN
                           => N741);
   U18713 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_16_port, A2 => n11814, ZN
                           => N742);
   U18714 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_17_port, A2 => n11814, ZN
                           => N743);
   U18715 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_18_port, A2 => n11814, ZN
                           => N744);
   U18716 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_19_port, A2 => n11814, ZN
                           => N745);
   U18717 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_20_port, A2 => n11814, ZN
                           => N746);
   U18718 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_21_port, A2 => n11814, ZN
                           => N747);
   U18719 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_22_port, A2 => n11814, ZN
                           => N748);
   U18720 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_23_port, A2 => n11814, ZN
                           => N749);
   U18721 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_24_port, A2 => n11814, ZN
                           => N750);
   U18722 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_25_port, A2 => n11814, ZN
                           => N751);
   U18723 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_26_port, A2 => n11815, ZN
                           => N752);
   U18724 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_27_port, A2 => n11815, ZN
                           => N753);
   U18725 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_28_port, A2 => n11815, ZN
                           => N754);
   U18726 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_29_port, A2 => n11815, ZN
                           => N755);
   U18727 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_30_port, A2 => n11815, ZN
                           => N756);
   U18728 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_31_port, A2 => n11815, ZN
                           => N757);
   U18729 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_32_port, A2 => n11815, ZN
                           => N758);
   U18730 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_33_port, A2 => n11815, ZN
                           => N759);
   U18731 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_34_port, A2 => n11815, ZN
                           => N760);
   U18732 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_35_port, A2 => n11815, ZN
                           => N761);
   U18733 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_36_port, A2 => n11815, ZN
                           => N762);
   U18734 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_37_port, A2 => n11816, ZN
                           => N763);
   U18735 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_38_port, A2 => n11816, ZN
                           => N764);
   U18736 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_39_port, A2 => n11816, ZN
                           => N765);
   U18737 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_40_port, A2 => n11816, ZN
                           => N766);
   U18738 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_41_port, A2 => n11816, ZN
                           => N767);
   U18739 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_42_port, A2 => n11816, ZN
                           => N768);
   U18740 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_43_port, A2 => n11816, ZN
                           => N769);
   U18741 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_44_port, A2 => n11816, ZN
                           => N770);
   U18742 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_45_port, A2 => n11816, ZN
                           => N771);
   U18743 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_46_port, A2 => n11816, ZN
                           => N772);
   U18744 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_47_port, A2 => n11816, ZN
                           => N773);
   U18745 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_48_port, A2 => n11817, ZN
                           => N774);
   U18746 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_49_port, A2 => n11817, ZN
                           => N775);
   U18747 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_50_port, A2 => n11817, ZN
                           => N776);
   U18748 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_51_port, A2 => n11817, ZN
                           => N777);
   U18749 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_52_port, A2 => n11817, ZN
                           => N778);
   U18750 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_53_port, A2 => n11817, ZN
                           => N779);
   U18751 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_54_port, A2 => n11817, ZN
                           => N780);
   U18752 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_55_port, A2 => n11817, ZN
                           => N781);
   U18753 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_56_port, A2 => n11817, ZN
                           => N782);
   U18754 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_57_port, A2 => n11817, ZN
                           => N783);
   U18755 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_58_port, A2 => n11817, ZN
                           => N784);
   U18756 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_59_port, A2 => n11818, ZN
                           => N785);
   U18757 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_60_port, A2 => n11818, ZN
                           => N786);
   U18758 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_61_port, A2 => n11818, ZN
                           => N787);
   U18759 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_62_port, A2 => n11818, ZN
                           => N788);
   U18760 : AND2_X1 port map( A1 => NEXT_REGISTERS_20_63_port, A2 => n11818, ZN
                           => N789);
   U18761 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_0_port, A2 => n11818, ZN 
                           => N790);
   U18762 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_1_port, A2 => n11818, ZN 
                           => N791);
   U18763 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_2_port, A2 => n11818, ZN 
                           => N792);
   U18764 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_3_port, A2 => n11818, ZN 
                           => N793);
   U18765 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_4_port, A2 => n11818, ZN 
                           => N794);
   U18766 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_5_port, A2 => n11818, ZN 
                           => N795);
   U18767 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_6_port, A2 => n11819, ZN 
                           => N796);
   U18768 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_7_port, A2 => n11819, ZN 
                           => N797);
   U18769 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_8_port, A2 => n11819, ZN 
                           => N798);
   U18770 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_9_port, A2 => n11819, ZN 
                           => N799);
   U18771 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_10_port, A2 => n11819, ZN
                           => N800);
   U18772 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_11_port, A2 => n11819, ZN
                           => N801);
   U18773 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_12_port, A2 => n11819, ZN
                           => N802);
   U18774 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_13_port, A2 => n11819, ZN
                           => N803);
   U18775 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_14_port, A2 => n11819, ZN
                           => N804);
   U18776 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_15_port, A2 => n11819, ZN
                           => N805);
   U18777 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_16_port, A2 => n11819, ZN
                           => N806);
   U18778 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_17_port, A2 => n11820, ZN
                           => N807);
   U18779 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_18_port, A2 => n11820, ZN
                           => N808);
   U18780 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_19_port, A2 => n11820, ZN
                           => N809);
   U18781 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_20_port, A2 => n11820, ZN
                           => N810);
   U18782 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_21_port, A2 => n11820, ZN
                           => N811);
   U18783 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_22_port, A2 => n11820, ZN
                           => N812);
   U18784 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_23_port, A2 => n11820, ZN
                           => N813);
   U18785 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_24_port, A2 => n11820, ZN
                           => N814);
   U18786 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_25_port, A2 => n11820, ZN
                           => N815);
   U18787 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_26_port, A2 => n11820, ZN
                           => N816);
   U18788 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_27_port, A2 => n11820, ZN
                           => N817);
   U18789 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_28_port, A2 => n11821, ZN
                           => N818);
   U18790 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_29_port, A2 => n11821, ZN
                           => N819);
   U18791 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_30_port, A2 => n11821, ZN
                           => N820);
   U18792 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_31_port, A2 => n11821, ZN
                           => N821);
   U18793 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_32_port, A2 => n11821, ZN
                           => N822);
   U18794 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_33_port, A2 => n11821, ZN
                           => N823);
   U18795 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_34_port, A2 => n11821, ZN
                           => N824);
   U18796 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_35_port, A2 => n11821, ZN
                           => N825);
   U18797 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_36_port, A2 => n11821, ZN
                           => N826);
   U18798 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_37_port, A2 => n11821, ZN
                           => N827);
   U18799 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_38_port, A2 => n11821, ZN
                           => N828);
   U18800 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_39_port, A2 => n11822, ZN
                           => N829);
   U18801 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_40_port, A2 => n11822, ZN
                           => N830);
   U18802 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_41_port, A2 => n11822, ZN
                           => N831);
   U18803 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_42_port, A2 => n11822, ZN
                           => N832);
   U18804 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_43_port, A2 => n11822, ZN
                           => N833);
   U18805 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_44_port, A2 => n11822, ZN
                           => N834);
   U18806 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_45_port, A2 => n11822, ZN
                           => N835);
   U18807 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_46_port, A2 => n11822, ZN
                           => N836);
   U18808 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_47_port, A2 => n11822, ZN
                           => N837);
   U18809 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_48_port, A2 => n11822, ZN
                           => N838);
   U18810 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_49_port, A2 => n11822, ZN
                           => N839);
   U18811 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_50_port, A2 => n11823, ZN
                           => N840);
   U18812 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_51_port, A2 => n11823, ZN
                           => N841);
   U18813 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_52_port, A2 => n11823, ZN
                           => N842);
   U18814 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_53_port, A2 => n11823, ZN
                           => N843);
   U18815 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_54_port, A2 => n11823, ZN
                           => N844);
   U18816 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_55_port, A2 => n11823, ZN
                           => N845);
   U18817 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_56_port, A2 => n11823, ZN
                           => N846);
   U18818 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_57_port, A2 => n11823, ZN
                           => N847);
   U18819 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_58_port, A2 => n11823, ZN
                           => N848);
   U18820 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_59_port, A2 => n11823, ZN
                           => N849);
   U18821 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_60_port, A2 => n11824, ZN
                           => N850);
   U18822 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_61_port, A2 => n11824, ZN
                           => N851);
   U18823 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_62_port, A2 => n11824, ZN
                           => N852);
   U18824 : AND2_X1 port map( A1 => NEXT_REGISTERS_19_63_port, A2 => n11824, ZN
                           => N853);
   U18825 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_0_port, A2 => n11824, ZN 
                           => N854);
   U18826 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_1_port, A2 => n11824, ZN 
                           => N855);
   U18827 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_2_port, A2 => n11824, ZN 
                           => N856);
   U18828 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_3_port, A2 => n11824, ZN 
                           => N857);
   U18829 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_4_port, A2 => n11824, ZN 
                           => N858);
   U18830 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_5_port, A2 => n11824, ZN 
                           => N859);
   U18831 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_6_port, A2 => n11824, ZN 
                           => N860);
   U18832 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_7_port, A2 => n11825, ZN 
                           => N861);
   U18833 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_8_port, A2 => n11825, ZN 
                           => N862);
   U18834 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_9_port, A2 => n11825, ZN 
                           => N863);
   U18835 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_10_port, A2 => n11825, ZN
                           => N864);
   U18836 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_11_port, A2 => n11825, ZN
                           => N865);
   U18837 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_12_port, A2 => n11825, ZN
                           => N866);
   U18838 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_13_port, A2 => n11825, ZN
                           => N867);
   U18839 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_14_port, A2 => n11825, ZN
                           => N868);
   U18840 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_15_port, A2 => n11825, ZN
                           => N869);
   U18841 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_16_port, A2 => n11825, ZN
                           => N870);
   U18842 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_17_port, A2 => n11825, ZN
                           => N871);
   U18843 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_18_port, A2 => n11826, ZN
                           => N872);
   U18844 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_19_port, A2 => n11826, ZN
                           => N873);
   U18845 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_20_port, A2 => n11826, ZN
                           => N874);
   U18846 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_21_port, A2 => n11826, ZN
                           => N875);
   U18847 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_22_port, A2 => n11826, ZN
                           => N876);
   U18848 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_23_port, A2 => n11826, ZN
                           => N877);
   U18849 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_24_port, A2 => n11826, ZN
                           => N878);
   U18850 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_25_port, A2 => n11826, ZN
                           => N879);
   U18851 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_26_port, A2 => n11826, ZN
                           => N880);
   U18852 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_27_port, A2 => n11826, ZN
                           => N881);
   U18853 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_28_port, A2 => n11826, ZN
                           => N882);
   U18854 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_29_port, A2 => n11827, ZN
                           => N883);
   U18855 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_30_port, A2 => n11827, ZN
                           => N884);
   U18856 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_31_port, A2 => n11827, ZN
                           => N885);
   U18857 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_32_port, A2 => n11827, ZN
                           => N886);
   U18858 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_33_port, A2 => n11827, ZN
                           => N887);
   U18859 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_34_port, A2 => n11827, ZN
                           => N888);
   U18860 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_35_port, A2 => n11827, ZN
                           => N889);
   U18861 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_36_port, A2 => n11827, ZN
                           => N890);
   U18862 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_37_port, A2 => n11827, ZN
                           => N891);
   U18863 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_38_port, A2 => n11827, ZN
                           => N892);
   U18864 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_39_port, A2 => n11827, ZN
                           => N893);
   U18865 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_40_port, A2 => n11828, ZN
                           => N894);
   U18866 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_41_port, A2 => n11828, ZN
                           => N895);
   U18867 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_42_port, A2 => n11828, ZN
                           => N896);
   U18868 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_43_port, A2 => n11828, ZN
                           => N897);
   U18869 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_44_port, A2 => n11828, ZN
                           => N898);
   U18870 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_45_port, A2 => n11828, ZN
                           => N899);
   U18871 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_46_port, A2 => n11828, ZN
                           => N900);
   U18872 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_47_port, A2 => n11828, ZN
                           => N901);
   U18873 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_48_port, A2 => n11828, ZN
                           => N902);
   U18874 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_49_port, A2 => n11828, ZN
                           => N903);
   U18875 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_50_port, A2 => n11828, ZN
                           => N904);
   U18876 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_51_port, A2 => n11829, ZN
                           => N905);
   U18877 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_52_port, A2 => n11829, ZN
                           => N906);
   U18878 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_53_port, A2 => n11829, ZN
                           => N907);
   U18879 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_54_port, A2 => n11829, ZN
                           => N908);
   U18880 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_55_port, A2 => n11829, ZN
                           => N909);
   U18881 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_56_port, A2 => n11829, ZN
                           => N910);
   U18882 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_57_port, A2 => n11829, ZN
                           => N911);
   U18883 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_58_port, A2 => n11829, ZN
                           => N912);
   U18884 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_59_port, A2 => n11829, ZN
                           => N913);
   U18885 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_60_port, A2 => n11829, ZN
                           => N914);
   U18886 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_61_port, A2 => n11829, ZN
                           => N915);
   U18887 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_62_port, A2 => n11830, ZN
                           => N916);
   U18888 : AND2_X1 port map( A1 => NEXT_REGISTERS_18_63_port, A2 => n11830, ZN
                           => N917);
   U18889 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_0_port, A2 => n11830, ZN 
                           => N918);
   U18890 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_1_port, A2 => n11830, ZN 
                           => N919);
   U18891 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_2_port, A2 => n11830, ZN 
                           => N920);
   U18892 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_3_port, A2 => n11830, ZN 
                           => N921);
   U18893 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_4_port, A2 => n11830, ZN 
                           => N922);
   U18894 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_5_port, A2 => n11830, ZN 
                           => N923);
   U18895 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_6_port, A2 => n11830, ZN 
                           => N924);
   U18896 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_7_port, A2 => n11830, ZN 
                           => N925);
   U18897 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_8_port, A2 => n11830, ZN 
                           => N926);
   U18898 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_9_port, A2 => n11831, ZN 
                           => N927);
   U18899 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_10_port, A2 => n11831, ZN
                           => N928);
   U18900 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_11_port, A2 => n11831, ZN
                           => N929);
   U18901 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_12_port, A2 => n11831, ZN
                           => N930);
   U18902 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_13_port, A2 => n11831, ZN
                           => N931);
   U18903 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_14_port, A2 => n11831, ZN
                           => N932);
   U18904 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_15_port, A2 => n11831, ZN
                           => N933);
   U18905 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_16_port, A2 => n11831, ZN
                           => N934);
   U18906 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_17_port, A2 => n11831, ZN
                           => N935);
   U18907 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_18_port, A2 => n11831, ZN
                           => N936);
   U18908 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_19_port, A2 => n11831, ZN
                           => N937);
   U18909 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_20_port, A2 => n11832, ZN
                           => N938);
   U18910 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_21_port, A2 => n11832, ZN
                           => N939);
   U18911 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_22_port, A2 => n11832, ZN
                           => N940);
   U18912 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_23_port, A2 => n11832, ZN
                           => N941);
   U18913 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_24_port, A2 => n11832, ZN
                           => N942);
   U18914 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_25_port, A2 => n11832, ZN
                           => N943);
   U18915 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_26_port, A2 => n11832, ZN
                           => N944);
   U18916 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_27_port, A2 => n11832, ZN
                           => N945);
   U18917 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_28_port, A2 => n11832, ZN
                           => N946);
   U18918 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_29_port, A2 => n11832, ZN
                           => N947);
   U18919 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_30_port, A2 => n11832, ZN
                           => N948);
   U18920 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_31_port, A2 => n11833, ZN
                           => N949);
   U18921 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_32_port, A2 => n11833, ZN
                           => N950);
   U18922 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_33_port, A2 => n11833, ZN
                           => N951);
   U18923 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_34_port, A2 => n11833, ZN
                           => N952);
   U18924 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_35_port, A2 => n11833, ZN
                           => N953);
   U18925 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_36_port, A2 => n11833, ZN
                           => N954);
   U18926 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_37_port, A2 => n11833, ZN
                           => N955);
   U18927 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_38_port, A2 => n11833, ZN
                           => N956);
   U18928 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_39_port, A2 => n11833, ZN
                           => N957);
   U18929 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_40_port, A2 => n11833, ZN
                           => N958);
   U18930 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_41_port, A2 => n11833, ZN
                           => N959);
   U18931 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_42_port, A2 => n11834, ZN
                           => N960);
   U18932 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_43_port, A2 => n11834, ZN
                           => N961);
   U18933 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_44_port, A2 => n11834, ZN
                           => N962);
   U18934 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_45_port, A2 => n11834, ZN
                           => N963);
   U18935 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_46_port, A2 => n11834, ZN
                           => N964);
   U18936 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_47_port, A2 => n11834, ZN
                           => N965);
   U18937 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_48_port, A2 => n11834, ZN
                           => N966);
   U18938 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_49_port, A2 => n11834, ZN
                           => N967);
   U18939 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_50_port, A2 => n11834, ZN
                           => N968);
   U18940 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_51_port, A2 => n11834, ZN
                           => N969);
   U18941 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_52_port, A2 => n11835, ZN
                           => N970);
   U18942 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_53_port, A2 => n11835, ZN
                           => N971);
   U18943 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_54_port, A2 => n11835, ZN
                           => N972);
   U18944 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_55_port, A2 => n11835, ZN
                           => N973);
   U18945 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_56_port, A2 => n11835, ZN
                           => N974);
   U18946 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_57_port, A2 => n11835, ZN
                           => N975);
   U18947 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_58_port, A2 => n11835, ZN
                           => N976);
   U18948 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_59_port, A2 => n11835, ZN
                           => N977);
   U18949 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_60_port, A2 => n11835, ZN
                           => N978);
   U18950 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_61_port, A2 => n11835, ZN
                           => N979);
   U18951 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_62_port, A2 => n11835, ZN
                           => N980);
   U18952 : AND2_X1 port map( A1 => NEXT_REGISTERS_17_63_port, A2 => n11836, ZN
                           => N981);
   U18953 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_0_port, A2 => n11836, ZN 
                           => N982);
   U18954 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_1_port, A2 => n11836, ZN 
                           => N983);
   U18955 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_2_port, A2 => n11836, ZN 
                           => N984);
   U18956 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_3_port, A2 => n11836, ZN 
                           => N985);
   U18957 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_4_port, A2 => n11836, ZN 
                           => N986);
   U18958 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_5_port, A2 => n11836, ZN 
                           => N987);
   U18959 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_6_port, A2 => n11836, ZN 
                           => N988);
   U18960 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_7_port, A2 => n11836, ZN 
                           => N989);
   U18961 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_8_port, A2 => n11836, ZN 
                           => N990);
   U18962 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_9_port, A2 => n11836, ZN 
                           => N991);
   U18963 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_10_port, A2 => n11837, ZN
                           => N992);
   U18964 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_11_port, A2 => n11837, ZN
                           => N993);
   U18965 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_12_port, A2 => n11837, ZN
                           => N994);
   U18966 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_13_port, A2 => n11837, ZN
                           => N995);
   U18967 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_14_port, A2 => n11837, ZN
                           => N996);
   U18968 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_15_port, A2 => n11837, ZN
                           => N997);
   U18969 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_16_port, A2 => n11837, ZN
                           => N998);
   U18970 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_17_port, A2 => n11837, ZN
                           => N999);
   U18971 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_18_port, A2 => n11667, ZN
                           => N1000);
   U18972 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_19_port, A2 => n11667, ZN
                           => N1001);
   U18973 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_20_port, A2 => n11667, ZN
                           => N1002);
   U18974 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_21_port, A2 => n11667, ZN
                           => N1003);
   U18975 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_22_port, A2 => n11667, ZN
                           => N1004);
   U18976 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_23_port, A2 => n11667, ZN
                           => N1005);
   U18977 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_24_port, A2 => n11667, ZN
                           => N1006);
   U18978 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_25_port, A2 => n11667, ZN
                           => N1007);
   U18979 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_26_port, A2 => n11667, ZN
                           => N1008);
   U18980 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_27_port, A2 => n11667, ZN
                           => N1009);
   U18981 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_28_port, A2 => n11668, ZN
                           => N1010);
   U18982 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_29_port, A2 => n11668, ZN
                           => N1011);
   U18983 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_30_port, A2 => n11668, ZN
                           => N1012);
   U18984 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_31_port, A2 => n11668, ZN
                           => N1013);
   U18985 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_32_port, A2 => n11668, ZN
                           => N1014);
   U18986 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_33_port, A2 => n11668, ZN
                           => N1015);
   U18987 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_34_port, A2 => n11668, ZN
                           => N1016);
   U18988 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_35_port, A2 => n11668, ZN
                           => N1017);
   U18989 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_36_port, A2 => n11668, ZN
                           => N1018);
   U18990 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_37_port, A2 => n11668, ZN
                           => N1019);
   U18991 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_38_port, A2 => n11668, ZN
                           => N1020);
   U18992 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_39_port, A2 => n11669, ZN
                           => N1021);
   U18993 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_40_port, A2 => n11669, ZN
                           => N1022);
   U18994 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_41_port, A2 => n11669, ZN
                           => N1023);
   U18995 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_42_port, A2 => n11669, ZN
                           => N1024);
   U18996 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_43_port, A2 => n11669, ZN
                           => N1025);
   U18997 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_44_port, A2 => n11669, ZN
                           => N1026);
   U18998 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_45_port, A2 => n11669, ZN
                           => N1027);
   U18999 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_46_port, A2 => n11669, ZN
                           => N1028);
   U19000 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_47_port, A2 => n11669, ZN
                           => N1029);
   U19001 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_48_port, A2 => n11669, ZN
                           => N1030);
   U19002 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_49_port, A2 => n11669, ZN
                           => N1031);
   U19003 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_50_port, A2 => n11670, ZN
                           => N1032);
   U19004 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_51_port, A2 => n11670, ZN
                           => N1033);
   U19005 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_52_port, A2 => n11670, ZN
                           => N1034);
   U19006 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_53_port, A2 => n11670, ZN
                           => N1035);
   U19007 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_54_port, A2 => n11670, ZN
                           => N1036);
   U19008 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_55_port, A2 => n11670, ZN
                           => N1037);
   U19009 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_56_port, A2 => n11670, ZN
                           => N1038);
   U19010 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_57_port, A2 => n11670, ZN
                           => N1039);
   U19011 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_58_port, A2 => n11670, ZN
                           => N1040);
   U19012 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_59_port, A2 => n11670, ZN
                           => N1041);
   U19013 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_60_port, A2 => n11670, ZN
                           => N1042);
   U19014 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_61_port, A2 => n11671, ZN
                           => N1043);
   U19015 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_62_port, A2 => n11671, ZN
                           => N1044);
   U19016 : AND2_X1 port map( A1 => NEXT_REGISTERS_16_63_port, A2 => n11671, ZN
                           => N1045);
   U19017 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_0_port, A2 => n11671, ZN 
                           => N1046);
   U19018 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_1_port, A2 => n11671, ZN 
                           => N1047);
   U19019 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_2_port, A2 => n11671, ZN 
                           => N1048);
   U19020 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_3_port, A2 => n11671, ZN 
                           => N1049);
   U19021 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_4_port, A2 => n11671, ZN 
                           => N1050);
   U19022 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_5_port, A2 => n11671, ZN 
                           => N1051);
   U19023 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_6_port, A2 => n11671, ZN 
                           => N1052);
   U19024 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_7_port, A2 => n11671, ZN 
                           => N1053);
   U19025 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_8_port, A2 => n11672, ZN 
                           => N1054);
   U19026 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_9_port, A2 => n11672, ZN 
                           => N1055);
   U19027 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_10_port, A2 => n11672, ZN
                           => N1056);
   U19028 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_11_port, A2 => n11672, ZN
                           => N1057);
   U19029 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_12_port, A2 => n11672, ZN
                           => N1058);
   U19030 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_13_port, A2 => n11672, ZN
                           => N1059);
   U19031 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_14_port, A2 => n11672, ZN
                           => N1060);
   U19032 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_15_port, A2 => n11672, ZN
                           => N1061);
   U19033 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_16_port, A2 => n11672, ZN
                           => N1062);
   U19034 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_17_port, A2 => n11672, ZN
                           => N1063);
   U19035 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_18_port, A2 => n11672, ZN
                           => N1064);
   U19036 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_19_port, A2 => n11673, ZN
                           => N1065);
   U19037 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_20_port, A2 => n11673, ZN
                           => N1066);
   U19038 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_21_port, A2 => n11673, ZN
                           => N1067);
   U19039 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_22_port, A2 => n11673, ZN
                           => N1068);
   U19040 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_23_port, A2 => n11673, ZN
                           => N1069);
   U19041 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_24_port, A2 => n11673, ZN
                           => N1070);
   U19042 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_25_port, A2 => n11673, ZN
                           => N1071);
   U19043 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_26_port, A2 => n11673, ZN
                           => N1072);
   U19044 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_27_port, A2 => n11673, ZN
                           => N1073);
   U19045 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_28_port, A2 => n11673, ZN
                           => N1074);
   U19046 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_29_port, A2 => n11673, ZN
                           => N1075);
   U19047 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_30_port, A2 => n11674, ZN
                           => N1076);
   U19048 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_31_port, A2 => n11674, ZN
                           => N1077);
   U19049 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_32_port, A2 => n11674, ZN
                           => N1078);
   U19050 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_33_port, A2 => n11674, ZN
                           => N1079);
   U19051 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_34_port, A2 => n11674, ZN
                           => N1080);
   U19052 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_35_port, A2 => n11674, ZN
                           => N1081);
   U19053 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_36_port, A2 => n11674, ZN
                           => N1082);
   U19054 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_37_port, A2 => n11674, ZN
                           => N1083);
   U19055 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_38_port, A2 => n11674, ZN
                           => N1084);
   U19056 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_39_port, A2 => n11674, ZN
                           => N1085);
   U19057 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_40_port, A2 => n11674, ZN
                           => N1086);
   U19058 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_41_port, A2 => n11675, ZN
                           => N1087);
   U19059 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_42_port, A2 => n11675, ZN
                           => N1088);
   U19060 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_43_port, A2 => n11675, ZN
                           => N1089);
   U19061 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_44_port, A2 => n11675, ZN
                           => N1090);
   U19062 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_45_port, A2 => n11675, ZN
                           => N1091);
   U19063 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_46_port, A2 => n11675, ZN
                           => N1092);
   U19064 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_47_port, A2 => n11675, ZN
                           => N1093);
   U19065 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_48_port, A2 => n11675, ZN
                           => N1094);
   U19066 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_49_port, A2 => n11675, ZN
                           => N1095);
   U19067 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_50_port, A2 => n11675, ZN
                           => N1096);
   U19068 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_51_port, A2 => n11675, ZN
                           => N1097);
   U19069 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_52_port, A2 => n11676, ZN
                           => N1098);
   U19070 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_53_port, A2 => n11676, ZN
                           => N1099);
   U19071 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_54_port, A2 => n11676, ZN
                           => N1100);
   U19072 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_55_port, A2 => n11676, ZN
                           => N1101);
   U19073 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_56_port, A2 => n11676, ZN
                           => N1102);
   U19074 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_57_port, A2 => n11676, ZN
                           => N1103);
   U19075 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_58_port, A2 => n11676, ZN
                           => N1104);
   U19076 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_59_port, A2 => n11676, ZN
                           => N1105);
   U19077 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_60_port, A2 => n11676, ZN
                           => N1106);
   U19078 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_61_port, A2 => n11676, ZN
                           => N1107);
   U19079 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_62_port, A2 => n11676, ZN
                           => N1108);
   U19080 : AND2_X1 port map( A1 => NEXT_REGISTERS_15_63_port, A2 => n11677, ZN
                           => N1109);
   U19081 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_0_port, A2 => n11677, ZN 
                           => N1110);
   U19082 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_1_port, A2 => n11677, ZN 
                           => N1111);
   U19083 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_2_port, A2 => n11677, ZN 
                           => N1112);
   U19084 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_3_port, A2 => n11677, ZN 
                           => N1113);
   U19085 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_4_port, A2 => n11677, ZN 
                           => N1114);
   U19086 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_5_port, A2 => n11677, ZN 
                           => N1115);
   U19087 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_6_port, A2 => n11677, ZN 
                           => N1116);
   U19088 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_7_port, A2 => n11677, ZN 
                           => N1117);
   U19089 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_8_port, A2 => n11677, ZN 
                           => N1118);
   U19090 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_9_port, A2 => n11677, ZN 
                           => N1119);
   U19091 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_10_port, A2 => n11678, ZN
                           => N1120);
   U19092 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_11_port, A2 => n11678, ZN
                           => N1121);
   U19093 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_12_port, A2 => n11678, ZN
                           => N1122);
   U19094 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_13_port, A2 => n11678, ZN
                           => N1123);
   U19095 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_14_port, A2 => n11678, ZN
                           => N1124);
   U19096 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_15_port, A2 => n11678, ZN
                           => N1125);
   U19097 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_16_port, A2 => n11678, ZN
                           => N1126);
   U19098 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_17_port, A2 => n11678, ZN
                           => N1127);
   U19099 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_18_port, A2 => n11678, ZN
                           => N1128);
   U19100 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_19_port, A2 => n11678, ZN
                           => N1129);
   U19101 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_20_port, A2 => n11679, ZN
                           => N1130);
   U19102 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_21_port, A2 => n11679, ZN
                           => N1131);
   U19103 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_22_port, A2 => n11679, ZN
                           => N1132);
   U19104 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_23_port, A2 => n11679, ZN
                           => N1133);
   U19105 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_24_port, A2 => n11679, ZN
                           => N1134);
   U19106 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_25_port, A2 => n11679, ZN
                           => N1135);
   U19107 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_26_port, A2 => n11679, ZN
                           => N1136);
   U19108 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_27_port, A2 => n11679, ZN
                           => N1137);
   U19109 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_28_port, A2 => n11679, ZN
                           => N1138);
   U19110 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_29_port, A2 => n11679, ZN
                           => N1139);
   U19111 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_30_port, A2 => n11679, ZN
                           => N1140);
   U19112 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_31_port, A2 => n11680, ZN
                           => N1141);
   U19113 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_32_port, A2 => n11680, ZN
                           => N1142);
   U19114 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_33_port, A2 => n11680, ZN
                           => N1143);
   U19115 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_34_port, A2 => n11680, ZN
                           => N1144);
   U19116 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_35_port, A2 => n11680, ZN
                           => N1145);
   U19117 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_36_port, A2 => n11680, ZN
                           => N1146);
   U19118 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_37_port, A2 => n11680, ZN
                           => N1147);
   U19119 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_38_port, A2 => n11680, ZN
                           => N1148);
   U19120 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_39_port, A2 => n11680, ZN
                           => N1149);
   U19121 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_40_port, A2 => n11680, ZN
                           => N1150);
   U19122 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_41_port, A2 => n11680, ZN
                           => N1151);
   U19123 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_42_port, A2 => n11681, ZN
                           => N1152);
   U19124 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_43_port, A2 => n11681, ZN
                           => N1153);
   U19125 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_44_port, A2 => n11681, ZN
                           => N1154);
   U19126 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_45_port, A2 => n11681, ZN
                           => N1155);
   U19127 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_46_port, A2 => n11681, ZN
                           => N1156);
   U19128 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_47_port, A2 => n11681, ZN
                           => N1157);
   U19129 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_48_port, A2 => n11681, ZN
                           => N1158);
   U19130 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_49_port, A2 => n11681, ZN
                           => N1159);
   U19131 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_50_port, A2 => n11681, ZN
                           => N1160);
   U19132 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_51_port, A2 => n11681, ZN
                           => N1161);
   U19133 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_52_port, A2 => n11681, ZN
                           => N1162);
   U19134 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_53_port, A2 => n11682, ZN
                           => N1163);
   U19135 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_54_port, A2 => n11682, ZN
                           => N1164);
   U19136 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_55_port, A2 => n11682, ZN
                           => N1165);
   U19137 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_56_port, A2 => n11682, ZN
                           => N1166);
   U19138 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_57_port, A2 => n11682, ZN
                           => N1167);
   U19139 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_58_port, A2 => n11682, ZN
                           => N1168);
   U19140 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_59_port, A2 => n11682, ZN
                           => N1169);
   U19141 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_60_port, A2 => n11682, ZN
                           => N1170);
   U19142 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_61_port, A2 => n11682, ZN
                           => N1171);
   U19143 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_62_port, A2 => n11682, ZN
                           => N1172);
   U19144 : AND2_X1 port map( A1 => NEXT_REGISTERS_14_63_port, A2 => n11682, ZN
                           => N1173);
   U19145 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_0_port, A2 => n11683, ZN 
                           => N1174);
   U19146 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_1_port, A2 => n11683, ZN 
                           => N1175);
   U19147 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_2_port, A2 => n11683, ZN 
                           => N1176);
   U19148 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_3_port, A2 => n11683, ZN 
                           => N1177);
   U19149 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_4_port, A2 => n11683, ZN 
                           => N1178);
   U19150 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_5_port, A2 => n11683, ZN 
                           => N1179);
   U19151 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_6_port, A2 => n11683, ZN 
                           => N1180);
   U19152 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_7_port, A2 => n11683, ZN 
                           => N1181);
   U19153 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_8_port, A2 => n11683, ZN 
                           => N1182);
   U19154 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_9_port, A2 => n11683, ZN 
                           => N1183);
   U19155 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_10_port, A2 => n11683, ZN
                           => N1184);
   U19156 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_11_port, A2 => n11684, ZN
                           => N1185);
   U19157 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_12_port, A2 => n11684, ZN
                           => N1186);
   U19158 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_13_port, A2 => n11684, ZN
                           => N1187);
   U19159 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_14_port, A2 => n11684, ZN
                           => N1188);
   U19160 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_15_port, A2 => n11684, ZN
                           => N1189);
   U19161 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_16_port, A2 => n11684, ZN
                           => N1190);
   U19162 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_17_port, A2 => n11684, ZN
                           => N1191);
   U19163 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_18_port, A2 => n11684, ZN
                           => N1192);
   U19164 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_19_port, A2 => n11684, ZN
                           => N1193);
   U19165 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_20_port, A2 => n11684, ZN
                           => N1194);
   U19166 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_21_port, A2 => n11684, ZN
                           => N1195);
   U19167 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_22_port, A2 => n11685, ZN
                           => N1196);
   U19168 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_23_port, A2 => n11685, ZN
                           => N1197);
   U19169 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_24_port, A2 => n11685, ZN
                           => N1198);
   U19170 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_25_port, A2 => n11685, ZN
                           => N1199);
   U19171 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_26_port, A2 => n11685, ZN
                           => N1200);
   U19172 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_27_port, A2 => n11685, ZN
                           => N1201);
   U19173 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_28_port, A2 => n11685, ZN
                           => N1202);
   U19174 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_29_port, A2 => n11685, ZN
                           => N1203);
   U19175 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_30_port, A2 => n11685, ZN
                           => N1204);
   U19176 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_31_port, A2 => n11685, ZN
                           => N1205);
   U19177 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_32_port, A2 => n11685, ZN
                           => N1206);
   U19178 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_33_port, A2 => n11686, ZN
                           => N1207);
   U19179 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_34_port, A2 => n11686, ZN
                           => N1208);
   U19180 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_35_port, A2 => n11686, ZN
                           => N1209);
   U19181 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_36_port, A2 => n11686, ZN
                           => N1210);
   U19182 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_37_port, A2 => n11686, ZN
                           => N1211);
   U19183 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_38_port, A2 => n11686, ZN
                           => N1212);
   U19184 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_39_port, A2 => n11686, ZN
                           => N1213);
   U19185 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_40_port, A2 => n11686, ZN
                           => N1214);
   U19186 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_41_port, A2 => n11686, ZN
                           => N1215);
   U19187 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_42_port, A2 => n11686, ZN
                           => N1216);
   U19188 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_43_port, A2 => n11686, ZN
                           => N1217);
   U19189 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_44_port, A2 => n11687, ZN
                           => N1218);
   U19190 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_45_port, A2 => n11687, ZN
                           => N1219);
   U19191 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_46_port, A2 => n11687, ZN
                           => N1220);
   U19192 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_47_port, A2 => n11687, ZN
                           => N1221);
   U19193 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_48_port, A2 => n11687, ZN
                           => N1222);
   U19194 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_49_port, A2 => n11687, ZN
                           => N1223);
   U19195 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_50_port, A2 => n11687, ZN
                           => N1224);
   U19196 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_51_port, A2 => n11687, ZN
                           => N1225);
   U19197 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_52_port, A2 => n11687, ZN
                           => N1226);
   U19198 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_53_port, A2 => n11687, ZN
                           => N1227);
   U19199 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_54_port, A2 => n11687, ZN
                           => N1228);
   U19200 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_55_port, A2 => n11688, ZN
                           => N1229);
   U19201 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_56_port, A2 => n11688, ZN
                           => N1230);
   U19202 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_57_port, A2 => n11688, ZN
                           => N1231);
   U19203 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_58_port, A2 => n11688, ZN
                           => N1232);
   U19204 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_59_port, A2 => n11688, ZN
                           => N1233);
   U19205 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_60_port, A2 => n11688, ZN
                           => N1234);
   U19206 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_61_port, A2 => n11688, ZN
                           => N1235);
   U19207 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_62_port, A2 => n11688, ZN
                           => N1236);
   U19208 : AND2_X1 port map( A1 => NEXT_REGISTERS_13_63_port, A2 => n11688, ZN
                           => N1237);
   U19209 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_0_port, A2 => n11688, ZN 
                           => N1238);
   U19210 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_1_port, A2 => n11688, ZN 
                           => N1239);
   U19211 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_2_port, A2 => n11689, ZN 
                           => N1240);
   U19212 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_3_port, A2 => n11689, ZN 
                           => N1241);
   U19213 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_4_port, A2 => n11689, ZN 
                           => N1242);
   U19214 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_5_port, A2 => n11689, ZN 
                           => N1243);
   U19215 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_6_port, A2 => n11689, ZN 
                           => N1244);
   U19216 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_7_port, A2 => n11689, ZN 
                           => N1245);
   U19217 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_8_port, A2 => n11689, ZN 
                           => N1246);
   U19218 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_9_port, A2 => n11689, ZN 
                           => N1247);
   U19219 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_10_port, A2 => n11689, ZN
                           => N1248);
   U19220 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_11_port, A2 => n11689, ZN
                           => N1249);
   U19221 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_12_port, A2 => n11690, ZN
                           => N1250);
   U19222 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_13_port, A2 => n11690, ZN
                           => N1251);
   U19223 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_14_port, A2 => n11690, ZN
                           => N1252);
   U19224 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_15_port, A2 => n11690, ZN
                           => N1253);
   U19225 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_16_port, A2 => n11690, ZN
                           => N1254);
   U19226 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_17_port, A2 => n11690, ZN
                           => N1255);
   U19227 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_18_port, A2 => n11690, ZN
                           => N1256);
   U19228 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_19_port, A2 => n11690, ZN
                           => N1257);
   U19229 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_20_port, A2 => n11690, ZN
                           => N1258);
   U19230 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_21_port, A2 => n11690, ZN
                           => N1259);
   U19231 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_22_port, A2 => n11690, ZN
                           => N1260);
   U19232 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_23_port, A2 => n11691, ZN
                           => N1261);
   U19233 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_24_port, A2 => n11691, ZN
                           => N1262);
   U19234 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_25_port, A2 => n11691, ZN
                           => N1263);
   U19235 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_26_port, A2 => n11691, ZN
                           => N1264);
   U19236 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_27_port, A2 => n11691, ZN
                           => N1265);
   U19237 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_28_port, A2 => n11691, ZN
                           => N1266);
   U19238 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_29_port, A2 => n11691, ZN
                           => N1267);
   U19239 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_30_port, A2 => n11691, ZN
                           => N1268);
   U19240 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_31_port, A2 => n11691, ZN
                           => N1269);
   U19241 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_32_port, A2 => n11691, ZN
                           => N1270);
   U19242 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_33_port, A2 => n11691, ZN
                           => N1271);
   U19243 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_34_port, A2 => n11692, ZN
                           => N1272);
   U19244 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_35_port, A2 => n11692, ZN
                           => N1273);
   U19245 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_36_port, A2 => n11692, ZN
                           => N1274);
   U19246 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_37_port, A2 => n11692, ZN
                           => N1275);
   U19247 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_38_port, A2 => n11692, ZN
                           => N1276);
   U19248 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_39_port, A2 => n11692, ZN
                           => N1277);
   U19249 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_40_port, A2 => n11692, ZN
                           => N1278);
   U19250 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_41_port, A2 => n11692, ZN
                           => N1279);
   U19251 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_42_port, A2 => n11692, ZN
                           => N1280);
   U19252 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_43_port, A2 => n11692, ZN
                           => N1281);
   U19253 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_44_port, A2 => n11692, ZN
                           => N1282);
   U19254 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_45_port, A2 => n11693, ZN
                           => N1283);
   U19255 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_46_port, A2 => n11693, ZN
                           => N1284);
   U19256 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_47_port, A2 => n11693, ZN
                           => N1285);
   U19257 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_48_port, A2 => n11693, ZN
                           => N1286);
   U19258 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_49_port, A2 => n11693, ZN
                           => N1287);
   U19259 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_50_port, A2 => n11693, ZN
                           => N1288);
   U19260 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_51_port, A2 => n11693, ZN
                           => N1289);
   U19261 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_52_port, A2 => n11693, ZN
                           => N1290);
   U19262 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_53_port, A2 => n11693, ZN
                           => N1291);
   U19263 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_54_port, A2 => n11693, ZN
                           => N1292);
   U19264 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_55_port, A2 => n11693, ZN
                           => N1293);
   U19265 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_56_port, A2 => n11694, ZN
                           => N1294);
   U19266 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_57_port, A2 => n11694, ZN
                           => N1295);
   U19267 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_58_port, A2 => n11694, ZN
                           => N1296);
   U19268 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_59_port, A2 => n11694, ZN
                           => N1297);
   U19269 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_60_port, A2 => n11694, ZN
                           => N1298);
   U19270 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_61_port, A2 => n11694, ZN
                           => N1299);
   U19271 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_62_port, A2 => n11694, ZN
                           => N1300);
   U19272 : AND2_X1 port map( A1 => NEXT_REGISTERS_12_63_port, A2 => n11694, ZN
                           => N1301);
   U19273 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_0_port, A2 => n11694, ZN 
                           => N1302);
   U19274 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_1_port, A2 => n11694, ZN 
                           => N1303);
   U19275 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_2_port, A2 => n11694, ZN 
                           => N1304);
   U19276 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_3_port, A2 => n11695, ZN 
                           => N1305);
   U19277 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_4_port, A2 => n11695, ZN 
                           => N1306);
   U19278 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_5_port, A2 => n11695, ZN 
                           => N1307);
   U19279 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_6_port, A2 => n11695, ZN 
                           => N1308);
   U19280 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_7_port, A2 => n11695, ZN 
                           => N1309);
   U19281 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_8_port, A2 => n11695, ZN 
                           => N1310);
   U19282 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_9_port, A2 => n11695, ZN 
                           => N1311);
   U19283 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_10_port, A2 => n11695, ZN
                           => N1312);
   U19284 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_11_port, A2 => n11695, ZN
                           => N1313);
   U19285 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_12_port, A2 => n11695, ZN
                           => N1314);
   U19286 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_13_port, A2 => n11695, ZN
                           => N1315);
   U19287 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_14_port, A2 => n11696, ZN
                           => N1316);
   U19288 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_15_port, A2 => n11696, ZN
                           => N1317);
   U19289 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_16_port, A2 => n11696, ZN
                           => N1318);
   U19290 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_17_port, A2 => n11696, ZN
                           => N1319);
   U19291 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_18_port, A2 => n11696, ZN
                           => N1320);
   U19292 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_19_port, A2 => n11696, ZN
                           => N1321);
   U19293 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_20_port, A2 => n11696, ZN
                           => N1322);
   U19294 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_21_port, A2 => n11696, ZN
                           => N1323);
   U19295 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_22_port, A2 => n11696, ZN
                           => N1324);
   U19296 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_23_port, A2 => n11696, ZN
                           => N1325);
   U19297 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_24_port, A2 => n11696, ZN
                           => N1326);
   U19298 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_25_port, A2 => n11697, ZN
                           => N1327);
   U19299 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_26_port, A2 => n11697, ZN
                           => N1328);
   U19300 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_27_port, A2 => n11697, ZN
                           => N1329);
   U19301 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_28_port, A2 => n11697, ZN
                           => N1330);
   U19302 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_29_port, A2 => n11697, ZN
                           => N1331);
   U19303 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_30_port, A2 => n11697, ZN
                           => N1332);
   U19304 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_31_port, A2 => n11697, ZN
                           => N1333);
   U19305 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_32_port, A2 => n11697, ZN
                           => N1334);
   U19306 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_33_port, A2 => n11697, ZN
                           => N1335);
   U19307 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_34_port, A2 => n11697, ZN
                           => N1336);
   U19308 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_35_port, A2 => n11697, ZN
                           => N1337);
   U19309 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_36_port, A2 => n11698, ZN
                           => N1338);
   U19310 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_37_port, A2 => n11698, ZN
                           => N1339);
   U19311 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_38_port, A2 => n11698, ZN
                           => N1340);
   U19312 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_39_port, A2 => n11698, ZN
                           => N1341);
   U19313 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_40_port, A2 => n11698, ZN
                           => N1342);
   U19314 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_41_port, A2 => n11698, ZN
                           => N1343);
   U19315 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_42_port, A2 => n11698, ZN
                           => N1344);
   U19316 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_43_port, A2 => n11698, ZN
                           => N1345);
   U19317 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_44_port, A2 => n11698, ZN
                           => N1346);
   U19318 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_45_port, A2 => n11698, ZN
                           => N1347);
   U19319 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_46_port, A2 => n11698, ZN
                           => N1348);
   U19320 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_47_port, A2 => n11699, ZN
                           => N1349);
   U19321 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_48_port, A2 => n11699, ZN
                           => N1350);
   U19322 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_49_port, A2 => n11699, ZN
                           => N1351);
   U19323 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_50_port, A2 => n11699, ZN
                           => N1352);
   U19324 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_51_port, A2 => n11699, ZN
                           => N1353);
   U19325 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_52_port, A2 => n11699, ZN
                           => N1354);
   U19326 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_53_port, A2 => n11699, ZN
                           => N1355);
   U19327 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_54_port, A2 => n11699, ZN
                           => N1356);
   U19328 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_55_port, A2 => n11699, ZN
                           => N1357);
   U19329 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_56_port, A2 => n11699, ZN
                           => N1358);
   U19330 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_57_port, A2 => n11699, ZN
                           => N1359);
   U19331 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_58_port, A2 => n11700, ZN
                           => N1360);
   U19332 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_59_port, A2 => n11700, ZN
                           => N1361);
   U19333 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_60_port, A2 => n11700, ZN
                           => N1362);
   U19334 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_61_port, A2 => n11700, ZN
                           => N1363);
   U19335 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_62_port, A2 => n11700, ZN
                           => N1364);
   U19336 : AND2_X1 port map( A1 => NEXT_REGISTERS_11_63_port, A2 => n11700, ZN
                           => N1365);
   U19337 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_0_port, A2 => n11700, ZN 
                           => N1366);
   U19338 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_1_port, A2 => n11700, ZN 
                           => N1367);
   U19339 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_2_port, A2 => n11700, ZN 
                           => N1368);
   U19340 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_3_port, A2 => n11700, ZN 
                           => N1369);
   U19341 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_4_port, A2 => n11701, ZN 
                           => N1370);
   U19342 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_5_port, A2 => n11701, ZN 
                           => N1371);
   U19343 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_6_port, A2 => n11701, ZN 
                           => N1372);
   U19344 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_7_port, A2 => n11701, ZN 
                           => N1373);
   U19345 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_8_port, A2 => n11701, ZN 
                           => N1374);
   U19346 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_9_port, A2 => n11701, ZN 
                           => N1375);
   U19347 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_10_port, A2 => n11701, ZN
                           => N1376);
   U19348 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_11_port, A2 => n11701, ZN
                           => N1377);
   U19349 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_12_port, A2 => n11701, ZN
                           => N1378);
   U19350 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_13_port, A2 => n11701, ZN
                           => N1379);
   U19351 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_14_port, A2 => n11701, ZN
                           => N1380);
   U19352 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_15_port, A2 => n11702, ZN
                           => N1381);
   U19353 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_16_port, A2 => n11702, ZN
                           => N1382);
   U19354 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_17_port, A2 => n11702, ZN
                           => N1383);
   U19355 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_18_port, A2 => n11702, ZN
                           => N1384);
   U19356 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_19_port, A2 => n11702, ZN
                           => N1385);
   U19357 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_20_port, A2 => n11702, ZN
                           => N1386);
   U19358 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_21_port, A2 => n11702, ZN
                           => N1387);
   U19359 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_22_port, A2 => n11702, ZN
                           => N1388);
   U19360 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_23_port, A2 => n11702, ZN
                           => N1389);
   U19361 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_24_port, A2 => n11702, ZN
                           => N1390);
   U19362 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_25_port, A2 => n11702, ZN
                           => N1391);
   U19363 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_26_port, A2 => n11703, ZN
                           => N1392);
   U19364 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_27_port, A2 => n11703, ZN
                           => N1393);
   U19365 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_28_port, A2 => n11703, ZN
                           => N1394);
   U19366 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_29_port, A2 => n11703, ZN
                           => N1395);
   U19367 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_30_port, A2 => n11703, ZN
                           => N1396);
   U19368 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_31_port, A2 => n11703, ZN
                           => N1397);
   U19369 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_32_port, A2 => n11703, ZN
                           => N1398);
   U19370 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_33_port, A2 => n11703, ZN
                           => N1399);
   U19371 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_34_port, A2 => n11703, ZN
                           => N1400);
   U19372 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_35_port, A2 => n11703, ZN
                           => N1401);
   U19373 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_36_port, A2 => n11703, ZN
                           => N1402);
   U19374 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_37_port, A2 => n11704, ZN
                           => N1403);
   U19375 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_38_port, A2 => n11704, ZN
                           => N1404);
   U19376 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_39_port, A2 => n11704, ZN
                           => N1405);
   U19377 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_40_port, A2 => n11704, ZN
                           => N1406);
   U19378 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_41_port, A2 => n11704, ZN
                           => N1407);
   U19379 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_42_port, A2 => n11704, ZN
                           => N1408);
   U19380 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_43_port, A2 => n11704, ZN
                           => N1409);
   U19381 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_44_port, A2 => n11704, ZN
                           => N1410);
   U19382 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_45_port, A2 => n11704, ZN
                           => N1411);
   U19383 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_46_port, A2 => n11704, ZN
                           => N1412);
   U19384 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_47_port, A2 => n11704, ZN
                           => N1413);
   U19385 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_48_port, A2 => n11705, ZN
                           => N1414);
   U19386 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_49_port, A2 => n11705, ZN
                           => N1415);
   U19387 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_50_port, A2 => n11705, ZN
                           => N1416);
   U19388 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_51_port, A2 => n11705, ZN
                           => N1417);
   U19389 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_52_port, A2 => n11705, ZN
                           => N1418);
   U19390 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_53_port, A2 => n11705, ZN
                           => N1419);
   U19391 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_54_port, A2 => n11705, ZN
                           => N1420);
   U19392 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_55_port, A2 => n11705, ZN
                           => N1421);
   U19393 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_56_port, A2 => n11705, ZN
                           => N1422);
   U19394 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_57_port, A2 => n11705, ZN
                           => N1423);
   U19395 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_58_port, A2 => n11705, ZN
                           => N1424);
   U19396 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_59_port, A2 => n11706, ZN
                           => N1425);
   U19397 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_60_port, A2 => n11706, ZN
                           => N1426);
   U19398 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_61_port, A2 => n11706, ZN
                           => N1427);
   U19399 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_62_port, A2 => n11706, ZN
                           => N1428);
   U19400 : AND2_X1 port map( A1 => NEXT_REGISTERS_10_63_port, A2 => n11706, ZN
                           => N1429);
   U19401 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_0_port, A2 => n11706, ZN 
                           => N1430);
   U19402 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_1_port, A2 => n11706, ZN 
                           => N1431);
   U19403 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_2_port, A2 => n11706, ZN 
                           => N1432);
   U19404 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_3_port, A2 => n11706, ZN 
                           => N1433);
   U19405 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_4_port, A2 => n11706, ZN 
                           => N1434);
   U19406 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_5_port, A2 => n11706, ZN 
                           => N1435);
   U19407 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_6_port, A2 => n11707, ZN 
                           => N1436);
   U19408 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_7_port, A2 => n11707, ZN 
                           => N1437);
   U19409 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_8_port, A2 => n11707, ZN 
                           => N1438);
   U19410 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_9_port, A2 => n11707, ZN 
                           => N1439);
   U19411 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_10_port, A2 => n11707, ZN 
                           => N1440);
   U19412 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_11_port, A2 => n11707, ZN 
                           => N1441);
   U19413 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_12_port, A2 => n11707, ZN 
                           => N1442);
   U19414 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_13_port, A2 => n11707, ZN 
                           => N1443);
   U19415 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_14_port, A2 => n11707, ZN 
                           => N1444);
   U19416 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_15_port, A2 => n11707, ZN 
                           => N1445);
   U19417 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_16_port, A2 => n11707, ZN 
                           => N1446);
   U19418 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_17_port, A2 => n11708, ZN 
                           => N1447);
   U19419 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_18_port, A2 => n11708, ZN 
                           => N1448);
   U19420 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_19_port, A2 => n11708, ZN 
                           => N1449);
   U19421 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_20_port, A2 => n11708, ZN 
                           => N1450);
   U19422 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_21_port, A2 => n11708, ZN 
                           => N1451);
   U19423 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_22_port, A2 => n11708, ZN 
                           => N1452);
   U19424 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_23_port, A2 => n11708, ZN 
                           => N1453);
   U19425 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_24_port, A2 => n11708, ZN 
                           => N1454);
   U19426 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_25_port, A2 => n11708, ZN 
                           => N1455);
   U19427 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_26_port, A2 => n11708, ZN 
                           => N1456);
   U19428 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_27_port, A2 => n11708, ZN 
                           => N1457);
   U19429 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_28_port, A2 => n11709, ZN 
                           => N1458);
   U19430 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_29_port, A2 => n11709, ZN 
                           => N1459);
   U19431 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_30_port, A2 => n11709, ZN 
                           => N1460);
   U19432 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_31_port, A2 => n11709, ZN 
                           => N1461);
   U19433 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_32_port, A2 => n11709, ZN 
                           => N1462);
   U19434 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_33_port, A2 => n11709, ZN 
                           => N1463);
   U19435 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_34_port, A2 => n11709, ZN 
                           => N1464);
   U19436 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_35_port, A2 => n11709, ZN 
                           => N1465);
   U19437 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_36_port, A2 => n11709, ZN 
                           => N1466);
   U19438 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_37_port, A2 => n11709, ZN 
                           => N1467);
   U19439 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_38_port, A2 => n11709, ZN 
                           => N1468);
   U19440 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_39_port, A2 => n11710, ZN 
                           => N1469);
   U19441 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_40_port, A2 => n11710, ZN 
                           => N1470);
   U19442 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_41_port, A2 => n11710, ZN 
                           => N1471);
   U19443 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_42_port, A2 => n11710, ZN 
                           => N1472);
   U19444 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_43_port, A2 => n11710, ZN 
                           => N1473);
   U19445 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_44_port, A2 => n11710, ZN 
                           => N1474);
   U19446 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_45_port, A2 => n11710, ZN 
                           => N1475);
   U19447 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_46_port, A2 => n11710, ZN 
                           => N1476);
   U19448 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_47_port, A2 => n11710, ZN 
                           => N1477);
   U19449 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_48_port, A2 => n11710, ZN 
                           => N1478);
   U19450 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_49_port, A2 => n11710, ZN 
                           => N1479);
   U19451 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_50_port, A2 => n11711, ZN 
                           => N1480);
   U19452 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_51_port, A2 => n11711, ZN 
                           => N1481);
   U19453 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_52_port, A2 => n11711, ZN 
                           => N1482);
   U19454 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_53_port, A2 => n11711, ZN 
                           => N1483);
   U19455 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_54_port, A2 => n11711, ZN 
                           => N1484);
   U19456 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_55_port, A2 => n11711, ZN 
                           => N1485);
   U19457 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_56_port, A2 => n11711, ZN 
                           => N1486);
   U19458 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_57_port, A2 => n11711, ZN 
                           => N1487);
   U19459 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_58_port, A2 => n11711, ZN 
                           => N1488);
   U19460 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_59_port, A2 => n11711, ZN 
                           => N1489);
   U19461 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_60_port, A2 => n11712, ZN 
                           => N1490);
   U19462 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_61_port, A2 => n11712, ZN 
                           => N1491);
   U19463 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_62_port, A2 => n11712, ZN 
                           => N1492);
   U19464 : AND2_X1 port map( A1 => NEXT_REGISTERS_9_63_port, A2 => n11712, ZN 
                           => N1493);
   U19465 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_0_port, A2 => n11712, ZN 
                           => N1494);
   U19466 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_1_port, A2 => n11712, ZN 
                           => N1495);
   U19467 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_2_port, A2 => n11712, ZN 
                           => N1496);
   U19468 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_3_port, A2 => n11712, ZN 
                           => N1497);
   U19469 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_4_port, A2 => n11712, ZN 
                           => N1498);
   U19470 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_5_port, A2 => n11712, ZN 
                           => N1499);
   U19471 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_6_port, A2 => n11712, ZN 
                           => N1500);
   U19472 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_7_port, A2 => n11713, ZN 
                           => N1501);
   U19473 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_8_port, A2 => n11713, ZN 
                           => N1502);
   U19474 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_9_port, A2 => n11713, ZN 
                           => N1503);
   U19475 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_10_port, A2 => n11713, ZN 
                           => N1504);
   U19476 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_11_port, A2 => n11713, ZN 
                           => N1505);
   U19477 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_12_port, A2 => n11713, ZN 
                           => N1506);
   U19478 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_13_port, A2 => n11713, ZN 
                           => N1507);
   U19479 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_14_port, A2 => n11713, ZN 
                           => N1508);
   U19480 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_15_port, A2 => n11713, ZN 
                           => N1509);
   U19481 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_16_port, A2 => n11713, ZN 
                           => N1510);
   U19482 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_17_port, A2 => n11713, ZN 
                           => N1511);
   U19483 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_18_port, A2 => n11714, ZN 
                           => N1512);
   U19484 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_19_port, A2 => n11714, ZN 
                           => N1513);
   U19485 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_20_port, A2 => n11714, ZN 
                           => N1514);
   U19486 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_21_port, A2 => n11714, ZN 
                           => N1515);
   U19487 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_22_port, A2 => n11714, ZN 
                           => N1516);
   U19488 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_23_port, A2 => n11714, ZN 
                           => N1517);
   U19489 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_24_port, A2 => n11714, ZN 
                           => N1518);
   U19490 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_25_port, A2 => n11714, ZN 
                           => N1519);
   U19491 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_26_port, A2 => n11714, ZN 
                           => N1520);
   U19492 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_27_port, A2 => n11714, ZN 
                           => N1521);
   U19493 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_28_port, A2 => n11714, ZN 
                           => N1522);
   U19494 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_29_port, A2 => n11715, ZN 
                           => N1523);
   U19495 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_30_port, A2 => n11715, ZN 
                           => N1524);
   U19496 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_31_port, A2 => n11715, ZN 
                           => N1525);
   U19497 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_32_port, A2 => n11715, ZN 
                           => N1526);
   U19498 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_33_port, A2 => n11715, ZN 
                           => N1527);
   U19499 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_34_port, A2 => n11715, ZN 
                           => N1528);
   U19500 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_35_port, A2 => n11715, ZN 
                           => N1529);
   U19501 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_36_port, A2 => n11715, ZN 
                           => N1530);
   U19502 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_37_port, A2 => n11715, ZN 
                           => N1531);
   U19503 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_38_port, A2 => n11715, ZN 
                           => N1532);
   U19504 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_39_port, A2 => n11715, ZN 
                           => N1533);
   U19505 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_40_port, A2 => n11716, ZN 
                           => N1534);
   U19506 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_41_port, A2 => n11716, ZN 
                           => N1535);
   U19507 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_42_port, A2 => n11716, ZN 
                           => N1536);
   U19508 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_43_port, A2 => n11716, ZN 
                           => N1537);
   U19509 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_44_port, A2 => n11716, ZN 
                           => N1538);
   U19510 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_45_port, A2 => n11716, ZN 
                           => N1539);
   U19511 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_46_port, A2 => n11716, ZN 
                           => N1540);
   U19512 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_47_port, A2 => n11716, ZN 
                           => N1541);
   U19513 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_48_port, A2 => n11716, ZN 
                           => N1542);
   U19514 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_49_port, A2 => n11716, ZN 
                           => N1543);
   U19515 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_50_port, A2 => n11716, ZN 
                           => N1544);
   U19516 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_51_port, A2 => n11717, ZN 
                           => N1545);
   U19517 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_52_port, A2 => n11717, ZN 
                           => N1546);
   U19518 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_53_port, A2 => n11717, ZN 
                           => N1547);
   U19519 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_54_port, A2 => n11717, ZN 
                           => N1548);
   U19520 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_55_port, A2 => n11717, ZN 
                           => N1549);
   U19521 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_56_port, A2 => n11717, ZN 
                           => N1550);
   U19522 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_57_port, A2 => n11717, ZN 
                           => N1551);
   U19523 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_58_port, A2 => n11717, ZN 
                           => N1552);
   U19524 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_59_port, A2 => n11717, ZN 
                           => N1553);
   U19525 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_60_port, A2 => n11717, ZN 
                           => N1554);
   U19526 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_61_port, A2 => n11717, ZN 
                           => N1555);
   U19527 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_62_port, A2 => n11718, ZN 
                           => N1556);
   U19528 : AND2_X1 port map( A1 => NEXT_REGISTERS_8_63_port, A2 => n11718, ZN 
                           => N1557);
   U19529 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_0_port, A2 => n11718, ZN 
                           => N1558);
   U19530 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_1_port, A2 => n11718, ZN 
                           => N1559);
   U19531 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_2_port, A2 => n11718, ZN 
                           => N1560);
   U19532 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_3_port, A2 => n11718, ZN 
                           => N1561);
   U19533 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_4_port, A2 => n11718, ZN 
                           => N1562);
   U19534 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_5_port, A2 => n11718, ZN 
                           => N1563);
   U19535 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_6_port, A2 => n11718, ZN 
                           => N1564);
   U19536 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_7_port, A2 => n11718, ZN 
                           => N1565);
   U19537 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_8_port, A2 => n11718, ZN 
                           => N1566);
   U19538 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_9_port, A2 => n11719, ZN 
                           => N1567);
   U19539 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_10_port, A2 => n11719, ZN 
                           => N1568);
   U19540 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_11_port, A2 => n11719, ZN 
                           => N1569);
   U19541 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_12_port, A2 => n11719, ZN 
                           => N1570);
   U19542 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_13_port, A2 => n11719, ZN 
                           => N1571);
   U19543 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_14_port, A2 => n11719, ZN 
                           => N1572);
   U19544 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_15_port, A2 => n11719, ZN 
                           => N1573);
   U19545 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_16_port, A2 => n11719, ZN 
                           => N1574);
   U19546 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_17_port, A2 => n11719, ZN 
                           => N1575);
   U19547 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_18_port, A2 => n11719, ZN 
                           => N1576);
   U19548 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_19_port, A2 => n11719, ZN 
                           => N1577);
   U19549 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_20_port, A2 => n11720, ZN 
                           => N1578);
   U19550 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_21_port, A2 => n11720, ZN 
                           => N1579);
   U19551 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_22_port, A2 => n11720, ZN 
                           => N1580);
   U19552 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_23_port, A2 => n11720, ZN 
                           => N1581);
   U19553 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_24_port, A2 => n11720, ZN 
                           => N1582);
   U19554 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_25_port, A2 => n11720, ZN 
                           => N1583);
   U19555 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_26_port, A2 => n11720, ZN 
                           => N1584);
   U19556 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_27_port, A2 => n11720, ZN 
                           => N1585);
   U19557 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_28_port, A2 => n11720, ZN 
                           => N1586);
   U19558 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_29_port, A2 => n11720, ZN 
                           => N1587);
   U19559 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_30_port, A2 => n11720, ZN 
                           => N1588);
   U19560 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_31_port, A2 => n11721, ZN 
                           => N1589);
   U19561 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_32_port, A2 => n11721, ZN 
                           => N1590);
   U19562 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_33_port, A2 => n11721, ZN 
                           => N1591);
   U19563 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_34_port, A2 => n11721, ZN 
                           => N1592);
   U19564 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_35_port, A2 => n11721, ZN 
                           => N1593);
   U19565 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_36_port, A2 => n11721, ZN 
                           => N1594);
   U19566 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_37_port, A2 => n11721, ZN 
                           => N1595);
   U19567 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_38_port, A2 => n11721, ZN 
                           => N1596);
   U19568 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_39_port, A2 => n11721, ZN 
                           => N1597);
   U19569 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_40_port, A2 => n11721, ZN 
                           => N1598);
   U19570 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_41_port, A2 => n11721, ZN 
                           => N1599);
   U19571 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_42_port, A2 => n11722, ZN 
                           => N1600);
   U19572 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_43_port, A2 => n11722, ZN 
                           => N1601);
   U19573 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_44_port, A2 => n11722, ZN 
                           => N1602);
   U19574 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_45_port, A2 => n11722, ZN 
                           => N1603);
   U19575 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_46_port, A2 => n11722, ZN 
                           => N1604);
   U19576 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_47_port, A2 => n11722, ZN 
                           => N1605);
   U19577 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_48_port, A2 => n11722, ZN 
                           => N1606);
   U19578 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_49_port, A2 => n11722, ZN 
                           => N1607);
   U19579 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_50_port, A2 => n11722, ZN 
                           => N1608);
   U19580 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_51_port, A2 => n11722, ZN 
                           => N1609);
   U19581 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_52_port, A2 => n11723, ZN 
                           => N1610);
   U19582 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_53_port, A2 => n11723, ZN 
                           => N1611);
   U19583 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_54_port, A2 => n11723, ZN 
                           => N1612);
   U19584 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_55_port, A2 => n11723, ZN 
                           => N1613);
   U19585 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_56_port, A2 => n11723, ZN 
                           => N1614);
   U19586 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_57_port, A2 => n11723, ZN 
                           => N1615);
   U19587 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_58_port, A2 => n11723, ZN 
                           => N1616);
   U19588 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_59_port, A2 => n11723, ZN 
                           => N1617);
   U19589 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_60_port, A2 => n11723, ZN 
                           => N1618);
   U19590 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_61_port, A2 => n11723, ZN 
                           => N1619);
   U19591 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_62_port, A2 => n11723, ZN 
                           => N1620);
   U19592 : AND2_X1 port map( A1 => NEXT_REGISTERS_7_63_port, A2 => n11724, ZN 
                           => N1621);
   U19593 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_0_port, A2 => n11724, ZN 
                           => N1622);
   U19594 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_1_port, A2 => n11724, ZN 
                           => N1623);
   U19595 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_2_port, A2 => n11724, ZN 
                           => N1624);
   U19596 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_3_port, A2 => n11724, ZN 
                           => N1625);
   U19597 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_4_port, A2 => n11724, ZN 
                           => N1626);
   U19598 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_5_port, A2 => n11724, ZN 
                           => N1627);
   U19599 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_6_port, A2 => n11724, ZN 
                           => N1628);
   U19600 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_7_port, A2 => n11724, ZN 
                           => N1629);
   U19601 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_8_port, A2 => n11724, ZN 
                           => N1630);
   U19602 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_9_port, A2 => n11724, ZN 
                           => N1631);
   U19603 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_10_port, A2 => n11725, ZN 
                           => N1632);
   U19604 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_11_port, A2 => n11725, ZN 
                           => N1633);
   U19605 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_12_port, A2 => n11725, ZN 
                           => N1634);
   U19606 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_13_port, A2 => n11725, ZN 
                           => N1635);
   U19607 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_14_port, A2 => n11725, ZN 
                           => N1636);
   U19608 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_15_port, A2 => n11725, ZN 
                           => N1637);
   U19609 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_16_port, A2 => n11725, ZN 
                           => N1638);
   U19610 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_17_port, A2 => n11725, ZN 
                           => N1639);
   U19611 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_18_port, A2 => n11725, ZN 
                           => N1640);
   U19612 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_19_port, A2 => n11725, ZN 
                           => N1641);
   U19613 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_20_port, A2 => n11725, ZN 
                           => N1642);
   U19614 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_21_port, A2 => n11726, ZN 
                           => N1643);
   U19615 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_22_port, A2 => n11726, ZN 
                           => N1644);
   U19616 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_23_port, A2 => n11726, ZN 
                           => N1645);
   U19617 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_24_port, A2 => n11726, ZN 
                           => N1646);
   U19618 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_25_port, A2 => n11726, ZN 
                           => N1647);
   U19619 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_26_port, A2 => n11726, ZN 
                           => N1648);
   U19620 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_27_port, A2 => n11726, ZN 
                           => N1649);
   U19621 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_28_port, A2 => n11726, ZN 
                           => N1650);
   U19622 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_29_port, A2 => n11726, ZN 
                           => N1651);
   U19623 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_30_port, A2 => n11726, ZN 
                           => N1652);
   U19624 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_31_port, A2 => n11726, ZN 
                           => N1653);
   U19625 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_32_port, A2 => n11727, ZN 
                           => N1654);
   U19626 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_33_port, A2 => n11727, ZN 
                           => N1655);
   U19627 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_34_port, A2 => n11727, ZN 
                           => N1656);
   U19628 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_35_port, A2 => n11727, ZN 
                           => N1657);
   U19629 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_36_port, A2 => n11727, ZN 
                           => N1658);
   U19630 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_37_port, A2 => n11727, ZN 
                           => N1659);
   U19631 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_38_port, A2 => n11727, ZN 
                           => N1660);
   U19632 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_39_port, A2 => n11727, ZN 
                           => N1661);
   U19633 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_40_port, A2 => n11727, ZN 
                           => N1662);
   U19634 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_41_port, A2 => n11727, ZN 
                           => N1663);
   U19635 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_42_port, A2 => n11727, ZN 
                           => N1664);
   U19636 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_43_port, A2 => n11728, ZN 
                           => N1665);
   U19637 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_44_port, A2 => n11728, ZN 
                           => N1666);
   U19638 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_45_port, A2 => n11728, ZN 
                           => N1667);
   U19639 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_46_port, A2 => n11728, ZN 
                           => N1668);
   U19640 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_47_port, A2 => n11728, ZN 
                           => N1669);
   U19641 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_48_port, A2 => n11728, ZN 
                           => N1670);
   U19642 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_49_port, A2 => n11728, ZN 
                           => N1671);
   U19643 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_50_port, A2 => n11728, ZN 
                           => N1672);
   U19644 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_51_port, A2 => n11728, ZN 
                           => N1673);
   U19645 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_52_port, A2 => n11728, ZN 
                           => N1674);
   U19646 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_53_port, A2 => n11728, ZN 
                           => N1675);
   U19647 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_54_port, A2 => n11729, ZN 
                           => N1676);
   U19648 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_55_port, A2 => n11729, ZN 
                           => N1677);
   U19649 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_56_port, A2 => n11729, ZN 
                           => N1678);
   U19650 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_57_port, A2 => n11729, ZN 
                           => N1679);
   U19651 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_58_port, A2 => n11729, ZN 
                           => N1680);
   U19652 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_59_port, A2 => n11729, ZN 
                           => N1681);
   U19653 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_60_port, A2 => n11729, ZN 
                           => N1682);
   U19654 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_61_port, A2 => n11729, ZN 
                           => N1683);
   U19655 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_62_port, A2 => n11729, ZN 
                           => N1684);
   U19656 : AND2_X1 port map( A1 => NEXT_REGISTERS_6_63_port, A2 => n11729, ZN 
                           => N1685);
   U19657 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_0_port, A2 => n11729, ZN 
                           => N1686);
   U19658 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_1_port, A2 => n11730, ZN 
                           => N1687);
   U19659 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_2_port, A2 => n11730, ZN 
                           => N1688);
   U19660 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_3_port, A2 => n11730, ZN 
                           => N1689);
   U19661 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_4_port, A2 => n11730, ZN 
                           => N1690);
   U19662 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_5_port, A2 => n11730, ZN 
                           => N1691);
   U19663 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_6_port, A2 => n11730, ZN 
                           => N1692);
   U19664 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_7_port, A2 => n11730, ZN 
                           => N1693);
   U19665 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_8_port, A2 => n11730, ZN 
                           => N1694);
   U19666 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_9_port, A2 => n11730, ZN 
                           => N1695);
   U19667 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_10_port, A2 => n11730, ZN 
                           => N1696);
   U19668 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_11_port, A2 => n11730, ZN 
                           => N1697);
   U19669 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_12_port, A2 => n11731, ZN 
                           => N1698);
   U19670 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_13_port, A2 => n11731, ZN 
                           => N1699);
   U19671 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_14_port, A2 => n11731, ZN 
                           => N1700);
   U19672 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_15_port, A2 => n11731, ZN 
                           => N1701);
   U19673 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_16_port, A2 => n11731, ZN 
                           => N1702);
   U19674 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_17_port, A2 => n11731, ZN 
                           => N1703);
   U19675 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_18_port, A2 => n11731, ZN 
                           => N1704);
   U19676 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_19_port, A2 => n11731, ZN 
                           => N1705);
   U19677 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_20_port, A2 => n11731, ZN 
                           => N1706);
   U19678 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_21_port, A2 => n11731, ZN 
                           => N1707);
   U19679 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_22_port, A2 => n11731, ZN 
                           => N1708);
   U19680 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_23_port, A2 => n11732, ZN 
                           => N1709);
   U19681 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_24_port, A2 => n11732, ZN 
                           => N1710);
   U19682 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_25_port, A2 => n11732, ZN 
                           => N1711);
   U19683 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_26_port, A2 => n11732, ZN 
                           => N1712);
   U19684 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_27_port, A2 => n11732, ZN 
                           => N1713);
   U19685 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_28_port, A2 => n11732, ZN 
                           => N1714);
   U19686 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_29_port, A2 => n11732, ZN 
                           => N1715);
   U19687 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_30_port, A2 => n11732, ZN 
                           => N1716);
   U19688 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_31_port, A2 => n11732, ZN 
                           => N1717);
   U19689 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_32_port, A2 => n11732, ZN 
                           => N1718);
   U19690 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_33_port, A2 => n11732, ZN 
                           => N1719);
   U19691 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_34_port, A2 => n11733, ZN 
                           => N1720);
   U19692 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_35_port, A2 => n11733, ZN 
                           => N1721);
   U19693 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_36_port, A2 => n11733, ZN 
                           => N1722);
   U19694 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_37_port, A2 => n11733, ZN 
                           => N1723);
   U19695 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_38_port, A2 => n11733, ZN 
                           => N1724);
   U19696 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_39_port, A2 => n11733, ZN 
                           => N1725);
   U19697 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_40_port, A2 => n11733, ZN 
                           => N1726);
   U19698 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_41_port, A2 => n11733, ZN 
                           => N1727);
   U19699 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_42_port, A2 => n11733, ZN 
                           => N1728);
   U19700 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_43_port, A2 => n11733, ZN 
                           => N1729);
   U19701 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_44_port, A2 => n11734, ZN 
                           => N1730);
   U19702 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_45_port, A2 => n11734, ZN 
                           => N1731);
   U19703 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_46_port, A2 => n11734, ZN 
                           => N1732);
   U19704 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_47_port, A2 => n11734, ZN 
                           => N1733);
   U19705 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_48_port, A2 => n11734, ZN 
                           => N1734);
   U19706 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_49_port, A2 => n11734, ZN 
                           => N1735);
   U19707 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_50_port, A2 => n11734, ZN 
                           => N1736);
   U19708 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_51_port, A2 => n11734, ZN 
                           => N1737);
   U19709 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_52_port, A2 => n11734, ZN 
                           => N1738);
   U19710 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_53_port, A2 => n11734, ZN 
                           => N1739);
   U19711 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_54_port, A2 => n11734, ZN 
                           => N1740);
   U19712 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_55_port, A2 => n11735, ZN 
                           => N1741);
   U19713 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_56_port, A2 => n11735, ZN 
                           => N1742);
   U19714 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_57_port, A2 => n11735, ZN 
                           => N1743);
   U19715 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_58_port, A2 => n11735, ZN 
                           => N1744);
   U19716 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_59_port, A2 => n11735, ZN 
                           => N1745);
   U19717 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_60_port, A2 => n11735, ZN 
                           => N1746);
   U19718 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_61_port, A2 => n11735, ZN 
                           => N1747);
   U19719 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_62_port, A2 => n11735, ZN 
                           => N1748);
   U19720 : AND2_X1 port map( A1 => NEXT_REGISTERS_5_63_port, A2 => n11735, ZN 
                           => N1749);
   U19721 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_0_port, A2 => n11735, ZN 
                           => N1750);
   U19722 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_1_port, A2 => n11735, ZN 
                           => N1751);
   U19723 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_2_port, A2 => n11736, ZN 
                           => N1752);
   U19724 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_3_port, A2 => n11736, ZN 
                           => N1753);
   U19725 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_4_port, A2 => n11736, ZN 
                           => N1754);
   U19726 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_5_port, A2 => n11736, ZN 
                           => N1755);
   U19727 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_6_port, A2 => n11736, ZN 
                           => N1756);
   U19728 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_7_port, A2 => n11736, ZN 
                           => N1757);
   U19729 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_8_port, A2 => n11736, ZN 
                           => N1758);
   U19730 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_9_port, A2 => n11736, ZN 
                           => N1759);
   U19731 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_10_port, A2 => n11736, ZN 
                           => N1760);
   U19732 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_11_port, A2 => n11736, ZN 
                           => N1761);
   U19733 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_12_port, A2 => n11736, ZN 
                           => N1762);
   U19734 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_13_port, A2 => n11737, ZN 
                           => N1763);
   U19735 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_14_port, A2 => n11737, ZN 
                           => N1764);
   U19736 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_15_port, A2 => n11737, ZN 
                           => N1765);
   U19737 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_16_port, A2 => n11737, ZN 
                           => N1766);
   U19738 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_17_port, A2 => n11737, ZN 
                           => N1767);
   U19739 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_18_port, A2 => n11737, ZN 
                           => N1768);
   U19740 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_19_port, A2 => n11737, ZN 
                           => N1769);
   U19741 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_20_port, A2 => n11737, ZN 
                           => N1770);
   U19742 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_21_port, A2 => n11737, ZN 
                           => N1771);
   U19743 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_22_port, A2 => n11737, ZN 
                           => N1772);
   U19744 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_23_port, A2 => n11737, ZN 
                           => N1773);
   U19745 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_24_port, A2 => n11738, ZN 
                           => N1774);
   U19746 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_25_port, A2 => n11738, ZN 
                           => N1775);
   U19747 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_26_port, A2 => n11738, ZN 
                           => N1776);
   U19748 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_27_port, A2 => n11738, ZN 
                           => N1777);
   U19749 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_28_port, A2 => n11738, ZN 
                           => N1778);
   U19750 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_29_port, A2 => n11738, ZN 
                           => N1779);
   U19751 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_30_port, A2 => n11738, ZN 
                           => N1780);
   U19752 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_31_port, A2 => n11738, ZN 
                           => N1781);
   U19753 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_32_port, A2 => n11738, ZN 
                           => N1782);
   U19754 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_33_port, A2 => n11738, ZN 
                           => N1783);
   U19755 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_34_port, A2 => n11738, ZN 
                           => N1784);
   U19756 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_35_port, A2 => n11739, ZN 
                           => N1785);
   U19757 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_36_port, A2 => n11739, ZN 
                           => N1786);
   U19758 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_37_port, A2 => n11739, ZN 
                           => N1787);
   U19759 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_38_port, A2 => n11739, ZN 
                           => N1788);
   U19760 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_39_port, A2 => n11739, ZN 
                           => N1789);
   U19761 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_40_port, A2 => n11739, ZN 
                           => N1790);
   U19762 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_41_port, A2 => n11739, ZN 
                           => N1791);
   U19763 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_42_port, A2 => n11739, ZN 
                           => N1792);
   U19764 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_43_port, A2 => n11739, ZN 
                           => N1793);
   U19765 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_44_port, A2 => n11739, ZN 
                           => N1794);
   U19766 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_45_port, A2 => n11739, ZN 
                           => N1795);
   U19767 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_46_port, A2 => n11740, ZN 
                           => N1796);
   U19768 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_47_port, A2 => n11740, ZN 
                           => N1797);
   U19769 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_48_port, A2 => n11740, ZN 
                           => N1798);
   U19770 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_49_port, A2 => n11740, ZN 
                           => N1799);
   U19771 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_50_port, A2 => n11740, ZN 
                           => N1800);
   U19772 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_51_port, A2 => n11740, ZN 
                           => N1801);
   U19773 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_52_port, A2 => n11740, ZN 
                           => N1802);
   U19774 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_53_port, A2 => n11740, ZN 
                           => N1803);
   U19775 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_54_port, A2 => n11740, ZN 
                           => N1804);
   U19776 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_55_port, A2 => n11740, ZN 
                           => N1805);
   U19777 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_56_port, A2 => n11740, ZN 
                           => N1806);
   U19778 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_57_port, A2 => n11741, ZN 
                           => N1807);
   U19779 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_58_port, A2 => n11741, ZN 
                           => N1808);
   U19780 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_59_port, A2 => n11741, ZN 
                           => N1809);
   U19781 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_60_port, A2 => n11741, ZN 
                           => N1810);
   U19782 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_61_port, A2 => n11741, ZN 
                           => N1811);
   U19783 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_62_port, A2 => n11741, ZN 
                           => N1812);
   U19784 : AND2_X1 port map( A1 => NEXT_REGISTERS_4_63_port, A2 => n11741, ZN 
                           => N1813);
   U19785 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_0_port, A2 => n11741, ZN 
                           => N1814);
   U19786 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_1_port, A2 => n11741, ZN 
                           => N1815);
   U19787 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_2_port, A2 => n11741, ZN 
                           => N1816);
   U19788 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_3_port, A2 => n11741, ZN 
                           => N1817);
   U19789 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_4_port, A2 => n11742, ZN 
                           => N1818);
   U19790 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_5_port, A2 => n11742, ZN 
                           => N1819);
   U19791 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_6_port, A2 => n11742, ZN 
                           => N1820);
   U19792 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_7_port, A2 => n11742, ZN 
                           => N1821);
   U19793 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_8_port, A2 => n11742, ZN 
                           => N1822);
   U19794 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_9_port, A2 => n11742, ZN 
                           => N1823);
   U19795 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_10_port, A2 => n11742, ZN 
                           => N1824);
   U19796 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_11_port, A2 => n11742, ZN 
                           => N1825);
   U19797 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_12_port, A2 => n11742, ZN 
                           => N1826);
   U19798 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_13_port, A2 => n11742, ZN 
                           => N1827);
   U19799 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_14_port, A2 => n11742, ZN 
                           => N1828);
   U19800 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_15_port, A2 => n11743, ZN 
                           => N1829);
   U19801 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_16_port, A2 => n11743, ZN 
                           => N1830);
   U19802 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_17_port, A2 => n11743, ZN 
                           => N1831);
   U19803 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_18_port, A2 => n11743, ZN 
                           => N1832);
   U19804 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_19_port, A2 => n11743, ZN 
                           => N1833);
   U19805 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_20_port, A2 => n11743, ZN 
                           => N1834);
   U19806 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_21_port, A2 => n11743, ZN 
                           => N1835);
   U19807 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_22_port, A2 => n11743, ZN 
                           => N1836);
   U19808 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_23_port, A2 => n11743, ZN 
                           => N1837);
   U19809 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_24_port, A2 => n11743, ZN 
                           => N1838);
   U19810 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_25_port, A2 => n11743, ZN 
                           => N1839);
   U19811 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_26_port, A2 => n11744, ZN 
                           => N1840);
   U19812 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_27_port, A2 => n11744, ZN 
                           => N1841);
   U19813 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_28_port, A2 => n11744, ZN 
                           => N1842);
   U19814 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_29_port, A2 => n11744, ZN 
                           => N1843);
   U19815 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_30_port, A2 => n11744, ZN 
                           => N1844);
   U19816 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_31_port, A2 => n11744, ZN 
                           => N1845);
   U19817 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_32_port, A2 => n11744, ZN 
                           => N1846);
   U19818 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_33_port, A2 => n11744, ZN 
                           => N1847);
   U19819 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_34_port, A2 => n11744, ZN 
                           => N1848);
   U19820 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_35_port, A2 => n11744, ZN 
                           => N1849);
   U19821 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_36_port, A2 => n11745, ZN 
                           => N1850);
   U19822 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_37_port, A2 => n11745, ZN 
                           => N1851);
   U19823 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_38_port, A2 => n11745, ZN 
                           => N1852);
   U19824 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_39_port, A2 => n11745, ZN 
                           => N1853);
   U19825 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_40_port, A2 => n11745, ZN 
                           => N1854);
   U19826 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_41_port, A2 => n11745, ZN 
                           => N1855);
   U19827 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_42_port, A2 => n11745, ZN 
                           => N1856);
   U19828 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_43_port, A2 => n11745, ZN 
                           => N1857);
   U19829 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_44_port, A2 => n11745, ZN 
                           => N1858);
   U19830 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_45_port, A2 => n11745, ZN 
                           => N1859);
   U19831 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_46_port, A2 => n11745, ZN 
                           => N1860);
   U19832 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_47_port, A2 => n11746, ZN 
                           => N1861);
   U19833 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_48_port, A2 => n11746, ZN 
                           => N1862);
   U19834 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_49_port, A2 => n11746, ZN 
                           => N1863);
   U19835 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_50_port, A2 => n11746, ZN 
                           => N1864);
   U19836 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_51_port, A2 => n11746, ZN 
                           => N1865);
   U19837 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_52_port, A2 => n11746, ZN 
                           => N1866);
   U19838 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_53_port, A2 => n11746, ZN 
                           => N1867);
   U19839 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_54_port, A2 => n11746, ZN 
                           => N1868);
   U19840 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_55_port, A2 => n11746, ZN 
                           => N1869);
   U19841 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_56_port, A2 => n11746, ZN 
                           => N1870);
   U19842 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_57_port, A2 => n11746, ZN 
                           => N1871);
   U19843 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_58_port, A2 => n11747, ZN 
                           => N1872);
   U19844 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_59_port, A2 => n11747, ZN 
                           => N1873);
   U19845 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_60_port, A2 => n11747, ZN 
                           => N1874);
   U19846 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_61_port, A2 => n11747, ZN 
                           => N1875);
   U19847 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_62_port, A2 => n11747, ZN 
                           => N1876);
   U19848 : AND2_X1 port map( A1 => NEXT_REGISTERS_3_63_port, A2 => n11747, ZN 
                           => N1877);
   U19849 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_0_port, A2 => n11747, ZN 
                           => N1878);
   U19850 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_1_port, A2 => n11747, ZN 
                           => N1879);
   U19851 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_2_port, A2 => n11747, ZN 
                           => N1880);
   U19852 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_3_port, A2 => n11747, ZN 
                           => N1881);
   U19853 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_4_port, A2 => n11747, ZN 
                           => N1882);
   U19854 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_5_port, A2 => n11748, ZN 
                           => N1883);
   U19855 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_6_port, A2 => n11748, ZN 
                           => N1884);
   U19856 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_7_port, A2 => n11748, ZN 
                           => N1885);
   U19857 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_8_port, A2 => n11748, ZN 
                           => N1886);
   U19858 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_9_port, A2 => n11748, ZN 
                           => N1887);
   U19859 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_10_port, A2 => n11748, ZN 
                           => N1888);
   U19860 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_11_port, A2 => n11748, ZN 
                           => N1889);
   U19861 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_12_port, A2 => n11748, ZN 
                           => N1890);
   U19862 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_13_port, A2 => n11748, ZN 
                           => N1891);
   U19863 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_14_port, A2 => n11748, ZN 
                           => N1892);
   U19864 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_15_port, A2 => n11748, ZN 
                           => N1893);
   U19865 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_16_port, A2 => n11749, ZN 
                           => N1894);
   U19866 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_17_port, A2 => n11749, ZN 
                           => N1895);
   U19867 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_18_port, A2 => n11749, ZN 
                           => N1896);
   U19868 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_19_port, A2 => n11749, ZN 
                           => N1897);
   U19869 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_20_port, A2 => n11749, ZN 
                           => N1898);
   U19870 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_21_port, A2 => n11749, ZN 
                           => N1899);
   U19871 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_22_port, A2 => n11749, ZN 
                           => N1900);
   U19872 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_23_port, A2 => n11749, ZN 
                           => N1901);
   U19873 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_24_port, A2 => n11749, ZN 
                           => N1902);
   U19874 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_25_port, A2 => n11749, ZN 
                           => N1903);
   U19875 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_26_port, A2 => n11749, ZN 
                           => N1904);
   U19876 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_27_port, A2 => n11750, ZN 
                           => N1905);
   U19877 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_28_port, A2 => n11750, ZN 
                           => N1906);
   U19878 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_29_port, A2 => n11750, ZN 
                           => N1907);
   U19879 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_30_port, A2 => n11750, ZN 
                           => N1908);
   U19880 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_31_port, A2 => n11750, ZN 
                           => N1909);
   U19881 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_32_port, A2 => n11750, ZN 
                           => N1910);
   U19882 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_33_port, A2 => n11750, ZN 
                           => N1911);
   U19883 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_34_port, A2 => n11750, ZN 
                           => N1912);
   U19884 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_35_port, A2 => n11750, ZN 
                           => N1913);
   U19885 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_36_port, A2 => n11750, ZN 
                           => N1914);
   U19886 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_37_port, A2 => n11750, ZN 
                           => N1915);
   U19887 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_38_port, A2 => n11751, ZN 
                           => N1916);
   U19888 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_39_port, A2 => n11751, ZN 
                           => N1917);
   U19889 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_40_port, A2 => n11751, ZN 
                           => N1918);
   U19890 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_41_port, A2 => n11751, ZN 
                           => N1919);
   U19891 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_42_port, A2 => n11751, ZN 
                           => N1920);
   U19892 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_43_port, A2 => n11751, ZN 
                           => N1921);
   U19893 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_44_port, A2 => n11751, ZN 
                           => N1922);
   U19894 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_45_port, A2 => n11751, ZN 
                           => N1923);
   U19895 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_46_port, A2 => n11751, ZN 
                           => N1924);
   U19896 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_47_port, A2 => n11751, ZN 
                           => N1925);
   U19897 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_48_port, A2 => n11751, ZN 
                           => N1926);
   U19898 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_49_port, A2 => n11752, ZN 
                           => N1927);
   U19899 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_50_port, A2 => n11752, ZN 
                           => N1928);
   U19900 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_51_port, A2 => n11752, ZN 
                           => N1929);
   U19901 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_52_port, A2 => n11752, ZN 
                           => N1930);
   U19902 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_53_port, A2 => n11752, ZN 
                           => N1931);
   U19903 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_54_port, A2 => n11752, ZN 
                           => N1932);
   U19904 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_55_port, A2 => n11752, ZN 
                           => N1933);
   U19905 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_56_port, A2 => n11752, ZN 
                           => N1934);
   U19906 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_57_port, A2 => n11752, ZN 
                           => N1935);
   U19907 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_58_port, A2 => n11752, ZN 
                           => N1936);
   U19908 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_59_port, A2 => n11752, ZN 
                           => N1937);
   U19909 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_60_port, A2 => n11753, ZN 
                           => N1938);
   U19910 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_61_port, A2 => n11753, ZN 
                           => N1939);
   U19911 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_62_port, A2 => n11753, ZN 
                           => N1940);
   U19912 : AND2_X1 port map( A1 => NEXT_REGISTERS_2_63_port, A2 => n11753, ZN 
                           => N1941);
   U19913 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_0_port, A2 => n11753, ZN 
                           => N1942);
   U19914 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_1_port, A2 => n11753, ZN 
                           => N1943);
   U19915 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_2_port, A2 => n11753, ZN 
                           => N1944);
   U19916 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_3_port, A2 => n11753, ZN 
                           => N1945);
   U19917 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_4_port, A2 => n11753, ZN 
                           => N1946);
   U19918 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_5_port, A2 => n11753, ZN 
                           => N1947);
   U19919 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_6_port, A2 => n11753, ZN 
                           => N1948);
   U19920 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_7_port, A2 => n11754, ZN 
                           => N1949);
   U19921 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_8_port, A2 => n11754, ZN 
                           => N1950);
   U19922 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_9_port, A2 => n11754, ZN 
                           => N1951);
   U19923 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_10_port, A2 => n11754, ZN 
                           => N1952);
   U19924 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_11_port, A2 => n11754, ZN 
                           => N1953);
   U19925 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_12_port, A2 => n11754, ZN 
                           => N1954);
   U19926 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_13_port, A2 => n11754, ZN 
                           => N1955);
   U19927 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_14_port, A2 => n11754, ZN 
                           => N1956);
   U19928 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_15_port, A2 => n11754, ZN 
                           => N1957);
   U19929 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_16_port, A2 => n11754, ZN 
                           => N1958);
   U19930 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_17_port, A2 => n11754, ZN 
                           => N1959);
   U19931 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_18_port, A2 => n11755, ZN 
                           => N1960);
   U19932 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_19_port, A2 => n11755, ZN 
                           => N1961);
   U19933 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_20_port, A2 => n11755, ZN 
                           => N1962);
   U19934 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_21_port, A2 => n11755, ZN 
                           => N1963);
   U19935 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_22_port, A2 => n11755, ZN 
                           => N1964);
   U19936 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_23_port, A2 => n11755, ZN 
                           => N1965);
   U19937 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_24_port, A2 => n11755, ZN 
                           => N1966);
   U19938 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_25_port, A2 => n11755, ZN 
                           => N1967);
   U19939 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_26_port, A2 => n11755, ZN 
                           => N1968);
   U19940 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_27_port, A2 => n11755, ZN 
                           => N1969);
   U19941 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_28_port, A2 => n11756, ZN 
                           => N1970);
   U19942 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_29_port, A2 => n11756, ZN 
                           => N1971);
   U19943 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_30_port, A2 => n11756, ZN 
                           => N1972);
   U19944 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_31_port, A2 => n11756, ZN 
                           => N1973);
   U19945 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_32_port, A2 => n11756, ZN 
                           => N1974);
   U19946 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_33_port, A2 => n11756, ZN 
                           => N1975);
   U19947 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_34_port, A2 => n11756, ZN 
                           => N1976);
   U19948 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_35_port, A2 => n11756, ZN 
                           => N1977);
   U19949 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_36_port, A2 => n11756, ZN 
                           => N1978);
   U19950 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_37_port, A2 => n11756, ZN 
                           => N1979);
   U19951 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_38_port, A2 => n11756, ZN 
                           => N1980);
   U19952 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_39_port, A2 => n11757, ZN 
                           => N1981);
   U19953 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_40_port, A2 => n11757, ZN 
                           => N1982);
   U19954 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_41_port, A2 => n11757, ZN 
                           => N1983);
   U19955 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_42_port, A2 => n11757, ZN 
                           => N1984);
   U19956 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_43_port, A2 => n11757, ZN 
                           => N1985);
   U19957 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_44_port, A2 => n11757, ZN 
                           => N1986);
   U19958 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_45_port, A2 => n11757, ZN 
                           => N1987);
   U19959 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_46_port, A2 => n11757, ZN 
                           => N1988);
   U19960 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_47_port, A2 => n11757, ZN 
                           => N1989);
   U19961 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_48_port, A2 => n11757, ZN 
                           => N1990);
   U19962 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_49_port, A2 => n11757, ZN 
                           => N1991);
   U19963 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_50_port, A2 => n11758, ZN 
                           => N1992);
   U19964 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_51_port, A2 => n11758, ZN 
                           => N1993);
   U19965 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_52_port, A2 => n11758, ZN 
                           => N1994);
   U19966 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_53_port, A2 => n11758, ZN 
                           => N1995);
   U19967 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_54_port, A2 => n11758, ZN 
                           => N1996);
   U19968 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_55_port, A2 => n11758, ZN 
                           => N1997);
   U19969 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_56_port, A2 => n11758, ZN 
                           => N1998);
   U19970 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_57_port, A2 => n11758, ZN 
                           => N1999);
   U19971 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_58_port, A2 => n11758, ZN 
                           => N2000);
   U19972 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_59_port, A2 => n11758, ZN 
                           => N2001);
   U19973 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_60_port, A2 => n11758, ZN 
                           => N2002);
   U19974 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_61_port, A2 => n11759, ZN 
                           => N2003);
   U19975 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_62_port, A2 => n11759, ZN 
                           => N2004);
   U19976 : AND2_X1 port map( A1 => NEXT_REGISTERS_1_63_port, A2 => n11759, ZN 
                           => N2005);
   U19977 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_0_port, A2 => n11759, ZN 
                           => N2006);
   U19978 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_1_port, A2 => n11759, ZN 
                           => N2007);
   U19979 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_2_port, A2 => n11759, ZN 
                           => N2008);
   U19980 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_3_port, A2 => n11759, ZN 
                           => N2009);
   U19981 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_4_port, A2 => n11759, ZN 
                           => N2010);
   U19982 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_5_port, A2 => n11759, ZN 
                           => N2011);
   U19983 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_6_port, A2 => n11759, ZN 
                           => N2012);
   U19984 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_7_port, A2 => n11759, ZN 
                           => N2013);
   U19985 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_8_port, A2 => n11760, ZN 
                           => N2014);
   U19986 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_9_port, A2 => n11760, ZN 
                           => N2015);
   U19987 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_10_port, A2 => n11760, ZN 
                           => N2016);
   U19988 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_11_port, A2 => n11760, ZN 
                           => N2017);
   U19989 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_12_port, A2 => n11760, ZN 
                           => N2018);
   U19990 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_13_port, A2 => n11760, ZN 
                           => N2019);
   U19991 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_14_port, A2 => n11760, ZN 
                           => N2020);
   U19992 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_15_port, A2 => n11760, ZN 
                           => N2021);
   U19993 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_16_port, A2 => n11760, ZN 
                           => N2022);
   U19994 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_17_port, A2 => n11760, ZN 
                           => N2023);
   U19995 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_18_port, A2 => n11760, ZN 
                           => N2024);
   U19996 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_19_port, A2 => n11761, ZN 
                           => N2025);
   U19997 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_20_port, A2 => n11761, ZN 
                           => N2026);
   U19998 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_21_port, A2 => n11761, ZN 
                           => N2027);
   U19999 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_22_port, A2 => n11761, ZN 
                           => N2028);
   U20000 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_23_port, A2 => n11761, ZN 
                           => N2029);
   U20001 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_24_port, A2 => n11761, ZN 
                           => N2030);
   U20002 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_25_port, A2 => n11761, ZN 
                           => N2031);
   U20003 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_26_port, A2 => n11761, ZN 
                           => N2032);
   U20004 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_27_port, A2 => n11761, ZN 
                           => N2033);
   U20005 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_28_port, A2 => n11761, ZN 
                           => N2034);
   U20006 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_29_port, A2 => n11761, ZN 
                           => N2035);
   U20007 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_30_port, A2 => n11762, ZN 
                           => N2036);
   U20008 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_31_port, A2 => n11762, ZN 
                           => N2037);
   U20009 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_32_port, A2 => n11762, ZN 
                           => N2038);
   U20010 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_33_port, A2 => n11762, ZN 
                           => N2039);
   U20011 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_34_port, A2 => n11762, ZN 
                           => N2040);
   U20012 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_35_port, A2 => n11762, ZN 
                           => N2041);
   U20013 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_36_port, A2 => n11762, ZN 
                           => N2042);
   U20014 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_37_port, A2 => n11762, ZN 
                           => N2043);
   U20015 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_38_port, A2 => n11762, ZN 
                           => N2044);
   U20016 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_39_port, A2 => n11762, ZN 
                           => N2045);
   U20017 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_40_port, A2 => n11762, ZN 
                           => N2046);
   U20018 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_41_port, A2 => n11763, ZN 
                           => N2047);
   U20019 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_42_port, A2 => n11763, ZN 
                           => N2048);
   U20020 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_43_port, A2 => n11763, ZN 
                           => N2049);
   U20021 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_44_port, A2 => n11763, ZN 
                           => N2050);
   U20022 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_45_port, A2 => n11763, ZN 
                           => N2051);
   U20023 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_46_port, A2 => n11763, ZN 
                           => N2052);
   U20024 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_47_port, A2 => n11763, ZN 
                           => N2053);
   U20025 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_48_port, A2 => n11763, ZN 
                           => N2054);
   U20026 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_49_port, A2 => n11763, ZN 
                           => N2055);
   U20027 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_50_port, A2 => n11763, ZN 
                           => N2056);
   U20028 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_51_port, A2 => n11763, ZN 
                           => N2057);
   U20029 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_52_port, A2 => n11764, ZN 
                           => N2058);
   U20030 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_53_port, A2 => n11764, ZN 
                           => N2059);
   U20031 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_54_port, A2 => n11764, ZN 
                           => N2060);
   U20032 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_55_port, A2 => n11764, ZN 
                           => N2061);
   U20033 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_56_port, A2 => n11764, ZN 
                           => N2062);
   U20034 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_57_port, A2 => n11764, ZN 
                           => N2063);
   U20035 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_58_port, A2 => n11764, ZN 
                           => N2064);
   U20036 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_59_port, A2 => n11764, ZN 
                           => N2065);
   U20037 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_60_port, A2 => n11764, ZN 
                           => N2066);
   U20038 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_61_port, A2 => n11764, ZN 
                           => N2067);
   U20039 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_62_port, A2 => n11764, ZN 
                           => N2068);
   U20040 : AND2_X1 port map( A1 => NEXT_REGISTERS_0_63_port, A2 => n11765, ZN 
                           => N2069);

end SYN_A;

library IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE work.constants.ALL;

ENTITY P4_ADDER IS
  PORT (
		A   : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
		B   : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
    SUM : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0)
  );
END ENTITY P4_ADDER;

ARCHITECTURE STRUCT OF P4_ADDER IS

  COMPONENT CARRY_GENERATOR IS
    -- Generics changed to NBIT_PER_BLOCK and NBLOCKS to match the other TBs. 
    GENERIC (
      NBIT_PER_BLOCK : INTEGER := CARRY_SELECT_NBIT;
      NBLOCKS : INTEGER := SUM_GENERATOR_NBLOCKS);
    PORT (
      A : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
      B : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
      Cin : IN STD_LOGIC;
      Co : OUT STD_LOGIC_VECTOR(NBLOCKS - 1 DOWNTO 0));
  END COMPONENT;

  COMPONENT SUM_GENERATOR IS
    GENERIC (
      NBIT_PER_BLOCK : INTEGER := CARRY_SELECT_NBIT;
      NBLOCKS : INTEGER := SUM_GENERATOR_NBLOCKS);
    PORT (
      A : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
      B : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
          -- TODO: USE AN ARRAY FOR CI
      CI : IN STD_LOGIC_VECTOR(NBLOCKS - 1 DOWNTO 0);
      S : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0));
  END COMPONENT;

  
  SIGNAL cg_out: std_logic_vector(NBLOCKS - 1 DOWNTO 0);
BEGIN
  
  -- using default values for generics
  carry_net: CARRY_GENERATOR
  PORT MAP (
    A => A,
    B => B,
           );
  
  -- using default values for generics
  sum_gen: SUM_GENERATOR
  PORT MAP (
    -- A => 
    -- B =>
    S => SUM
           );

END ARCHITECTURE STRUCT;

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.constants.ALL;

ENTITY PG_NETWORK IS
	GENERIC (
		NBIT_PER_BLOCK : INTEGER := CARRY_SELECT_NBIT;
		NBLOCKS : INTEGER := SUM_GENERATOR_NBLOCK);
	PORT (
		A : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS - 1 DOWNTO 0);
		Cin : IN STD_LOGIC;
		g : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS DOWNTO 0);
		p : OUT STD_LOGIC_VECTOR(NBIT_PER_BLOCK * NBLOCKS DOWNTO 0));
		-- The -1 is not needed in g and p since they add one bit for the Cin
		-- 	and shift the others one position to the left.
END PG_NETWORK;

ARCHITECTURE BEHAVIORAL OF PG_NETWORK IS
BEGIN

	g <= (A AND B) & Cin;
	p <= (A XOR B) & '0';

END BEHAVIORAL;
